MPQ    �    h�  h                                                                                 �gH=��ʳ�5���2h��2@&Vk_u��ԭ(��x��
&�m6r��{e���U�.R��z�3s�2����N� DkmA�Xt�&�QQ�\mV���!��%��ɏT��G8�,#^��r��0��W|ׂ
�rW��Y�Elh� ��Lɣ~�LW@��������C/Yz�t!�	��)0��ER�5�a5��5�Gꔍs,��^Yr���6J���C<��H��������1R�@_h��	�V���?�,(���Pֶ�t��n��L�'����.���o���j��Mr�§Zv���J��ݽ"_�h��y������mMyP	�V���|y0.�z��4cY����Z����f̌[�$�&���2V�ݕ�cZk�mR`������ݽϲ�N�)��%(:�~���A^�-�E��z�����hLn �X����sD;����ro�f�fQ������>~�Ԏ�|z>�/�\�Z��r��״M�K����}͐�􅏐(�	h�N�j��E;�չ�ڂ��:�F�E���Xw��#�˪5oJ'�>_|��ԔfqV�����饉4��82�c�J6��ӣB,'l[�/��3�h�X�@��hB3����W��xB���v��Ҷ(|gx����U�G*:h�Tܬ�י.�sNa���}�("u
�ė"C��da2�Wu��3=�߂�ɷ@��:�V��ڎ�H7?iCx3���;_DP�?�\�	�2��s,T�z�~�	"9d:UU	~��<$�<�5�} <���/�Ů��~Z��7V}�𽁧�5e��Am�lP�I���0�f��(%�����8�O�:�&g\S��$o��\�-���s�w��0����8���zN��2���i����H��j�}vΡc��(����2�>��T GNks ���D���r��7Z4��۶H��F}}AI$�(z���jk��:���<ۻ��9
w�\�����?�}��U��`�8 F�1~���4Y��p+�Ks����v����=�U��H�t����]���>Hl�5j,�b�^'���4�褡�e��u_����x�bz-G4-�5��f��G�V{�)�����#�<�N��]��i���Jf�x#���g�L�QD�?hB���Z�Kp��n�YK6k����|�x��#Pb�R�M�w��t���\L._�a��GЈ��R�T�W�?&N!d�Լ�S�>�y�qS�����wq|�K�2$Xt\S�g��uC<�%����P��C(&��*�/
�1-%y�������K�)�P�`	���5d/)���	<oOÔ��g("�Ip-ex���KM
�c��
�H�L"�?S���j�#;(�C) S�m����MQ���`y:��>5Qv�6�8h�r�V�I>x�0e���l,X��s	�!�@�=]�(k���{���P3$�ܢ��{!�B�Y �=؇G{�<�]��t�)�/�8Z2`�:)�N6�/�����<G�p�%�S���b��De/�������Ƀ�!��c]�[p��t�;��/0�l1�'�h��]؄x����
���e����G$CP��>f&��`�H�[xS����V�~��蝶��Ğ#���~�H�uT|�̻z����m�ԣ����3��٩�ʰ����	xÊ�$�=m��1}��3,kfJ^Z�;���uTj3쉏ؑ�^��u�v7���;v�)%�]c��/�T�@�Rs
j��S���C����{��V�M���`V�ub�5�P�ޱog��,^G>^ϼ�����Y-���g�X6��Pt��?)�N���D����O�,�V}*�B;(�wI�wO��S[Ύ���M`���8��9:̱��:�������-~�z�Įa8�pQ��fQ?`�h/`L��ꤘH|&gY3�4u����)�0���(\mA�O xS+'��z��8�Μq�0�-RFa�p6$��V� �wH˯����z�y7�$P�r|�u���o1*AM��X���[�R�^�Rxk4k.T'�����R"�C7B�lq���J��(��9YTHG���ɜ^��� M0���BA��`���]���TbI}�f!�	)Wy%g_��U�� ��\Oq���y�����*y��7p����!�˗�u+�]� `b��Y#6V����	ak�MW�g$8�'�!Գ��,�Zr��`7�/���H� �/��������z�~GQ�B@O��k.����q��N�Ěۯ�M6�`�^n��*v9&�G��hԯCjj���cn�=Ĭq��LBÆ�7��>1!�2|>dT�bz!�zk�ܼ���5��$��>¹���{p��,r�*?%I�����"Щ�gN}����"��(x?1Rw?|�F�d�7Wo�̗�^"=��Uꝭ$XR<�e�:B�XR.C���T����c�����0�p��HP�"J���c�v� |G��&�K&��*�����:�O���h�g\y�U�R6�	+itKa�݁���l}*�Gel��_�V[;�S��$�LHO_p ݢ�";�Ն�nq~nE�G���j�a��XN�s� �'7�����}4ۗŌ��r5�A��] �Z����鹟�P�Du7�����b�5d ��t�q�A�j�ﭱ��In�XT7��x�1n8֥0 Iڣ�q������e3��K�d��%XN�e�5*B��7����B[ڦ��<V6�&���:*���
-��(dҢ�b�䒒!��0�mC���:F���� {���N}��"�,< ���	O� O<R����U�������A�yK���sùZ���3�t�4�����'Y]-S�'���Hk��-u�{��S�����0�~�V9�����}▥��?@��Uk�t��r�et�ts;̿�#��Nj��E��O	���ޣ�`Z�*m5b��Ū��F.^�@y��۸E��+���̌Vf����y�vnqz̡��0�w%BL6�kJ�/qbg|Ѥ�z��_�s�wi��}�`)�X��Zz=&��©k����68���匐N���_.{.��l��7�2�kFEi`y՚B���$�5"��E:b�2|cY�o��\K%�嚕�{X�4|0�*=2�0\��S��������¦�a[h�IA��?7��(ly(D�R����%!G_Q,4m�ܺ�����,�e�T��G�s	#Y/rDE�0l�H� �
2�ӽZ�$Yϼ�h�_R�G�'~�a@�&�"
M�q���x��t��Q��)�5�E
Q�|TWҰ���o�w,'y���q����J��7���c(2�����1��@���ۜ4V���|΋Gs�U�Ͷ�p��c�L�2���/��6?O8��J���U\h!�$��������"�����͵�8ک�	�^m(w	S�{r�wm�.v���pctbb�ԥ��`E��{$fr��j��`�����4�~�������M �
���MW�$d����9�i��ݒ�<E��� ���9�nk.Ȩ�?;�q���xfgw�����F@v~����י�����\��Zkcr�&���駆�x�k�O�ǐ�Kh���j�C����վȔ�~F����TΕ��D����o�b�>:��|���/4�V�e'�V+�D�4��2@�hJ����K�_�[�{z�&��h��@��dB�z�����Ԕz�-8�{邶�rx�n��*NG�6�RTQB� � .�U�a�w}��Q=Yr
x,G"gd�d�W38F��
@O���%���#9Fi��xΠy�6f7���^P�	��wK������`,�B����]W9lU���������XZm<2Q�/a�����Z������l��g��<A�1�Pwoa��	f��t(ୂ��r��|�R���Տ�\��?��-�����W��Y�қ��B�uY�P2�[N�ڂ���7N�Pߎ}Q�?�?1((<>��l�>@_� �s)\��t��՛��"�u4#`h�C��!��x �C��Ou2��x��uA��y���'
ҺȬ�%��/��ؗU� h�B_ �,~�&J�S��+qmK���t��v�KW�xq�4�R�o�+�H�~�}Fl �j���9�H�#uҷ�"������aɠ�Gx���z�}n-�;ɡ�qء/�Vv�@����]��#�Ծ|��Nӏ���5$�LJ�f�?��<���D���B��Z�����E.��	�k�kD���xh�P�R`eFR衯��j�.Z���DDM��xo�o�3W�E�&��*d<��m��>ߡ�q�����w��Xo��2���t�Kagm�_C7�O���/PR��(A��* (��5�y��r�;;�FN(��pl`�1t��u�/�V���3E<�]u��l[#�BImme3I�fx���0
b�L]]?����s�j���(D�G n$r�]0��#Q��,`��9Tpv5�8#�իq[�b���% �gl�n��n�'!4j�=��_�CW?�V��ԯk$+V[w$��v��B�� >آڷ���~)	ua8�u�5��N�)2u��������.Hc��UD �O����t���(����*�O5�� ����c�"��C���?����z鲏��emݷ7���}�9�&�5��Sl[��˷�=�YX��#�AMM��p���Y�0��|;�z^I�������T�Ǡ�,��P��qt�I��$�z�o�N=H���l��ΚfE����[�05300��SY�^������2�Y�v�6��G��) T
p
R��j]`��KܟA�:{���ʨ��[��`q��bW�)+1��I��P>Yr��%�����գjg�A�6�|ctG�\��C/N�j���ѓ��(,G�*��B�v���w�SVR���w`u8��[:G�N���g9��nKu�B����p����=?��
��L���3�D&b�RY���uv@�X�&��\� O�>�+"5~z.�)8���#�$?P2�aQa>�tp�U�B�[��H�?߻69�+��T�O$���|����1�5�MH	\�;���I��-�64�.�'T����R}��ܥ�Λ�>K���M9�_�H�Zm��b�^) aœ�F������8T�&��a�-	��%"Ѵ-�ٲ}9����U�ɇ�V��-*����`����Fyiu�m�. �E���q6�������k�VE��P�v����,ny%��RNኹ����J��5l碋L义r��ɘ��(�3H��,���i���VrM�o�W�_�:v4�h�7�#G�C�4�J�ne�Ȭ��q�ꆁ�������yrdo��b�yzFR����飋�Bڙ��n>Cp�e�rn�%$�Z��l��DYNx��&+Ϩ�;.Z��w�jF��+�r�.�g8C^�#��w���Q<��u:���R	�T���c����c�+��rp�NHk�KJ�%C�>�|�;�u{�&ĕO��|�_Q��6��O2pCE\@��ԛ6��i��h�����h��
*Ա�l��_h�M;�3���H
*$ ���"���amq����������bX	 8�*'��-����4S䌁�m�DA�!�]ۃ����d�J���DA��7Qm=�:�b�� dk�����$0���	I??:X�/g�s��n�a�0�?�@�9d��@���'(d�g� /�%�5��F�RI�Dځa5w=[B�����:��*��9�)�Q�����y!��08�K��9JFr��uH�{�_}�ɂ �����)\<����A�[���tҜ��,\S�d;���S��:ӹô]�<�/kI��*��]0P]�D+�b���ІC9zY���6��S�!\�a��~^�����dcR��{ɚ���/�t��r+�O�������;�G�Щ2��l��-��{;T��VU5=4�� �r��ǳ^�o��G��� u+��oV�)4��C��nltZ��
~�2�6LQ��J�bB끤H�8�D�-s�<��I�/��X0��Z���v��#/�B��63u��>u������_���.���l�-���>�F@Ăy0U��\�$���"��:=�[|��SoUa�K �Ě�?X�ż0�ҏ2M���nT�Tmِ� �����=rph�e�� $�7Y�G?�D��Ŝ����Q�o~m��C�"���nB@��T���Gn�#T��r���0'�����
�k��5��Y
T�h�"�BM~DOL@��O�=^!ID��s�Ϟ�tW���Ȭ)��E�Qpԗ�_�+���JQ�,b&���i����JV�����~R)�N͕�L1�o�@�qy��O1VS��x�Ëb2�С������&�L(]���uMt 
!�K��CY"�]ۧ����U���/�"3��RA�S�Ϻ�Bm�Z	�X�s�r�,.j	��i�Qc�8c��m��w)���$�}��I�ٻ���S����P�c��x�k�E�]��-�������ᮐ0zŒ�k�Ev���[���z`nz��c�c�?;��hD�fBڬ�(�����E~�4}�2��ͥ"\&�TZ�0nr��n�ú��!�s�Ҫ:@��;�h	3j|��ϝ�1�N�/ F���ޯc�e�;@o@�>>��|V���!V�3���h���}4�-2��J���I��b��[��(���*hP�@
�B�#�s�w��f���%v o�ވ�xoP��Eg�G s{���T��4�� .�W|a8^�}aH_X]-
�b"���d׶�W���33Ղ`�\@
zv���_���Z]i���xi���1�~��P��6Ò%��x��d},ʪ���]c��H9��5U�������22��3�
<m��/�Z���ZG��̎L����+����:�A�sP����/fT�I(�����*���bƽ���\������^ß-=R����^�z���vl��rU����%26���)������s�},����c(��Ħ���>��� ���sD����㬞�j.�]l�4�Qm�>5������ �^��ʟ����s��kߵտ����
-���g��b��sN?U�%���� |f�~��U�mL���SK�����tv�F��<��,5�jrT��ȷ�8 �l�j"����
�^K��B���+ҳ�A÷x��z#Դ-za$�ܳ��<8�Vq�s�@�+��#�i�8�N�`c�"Y�罷f�&)�R#�zD౱B��qZo#ߜ==���k��2ږx#��P7��Rۜ-Aǡꉦ��\.U|�Ɵ`ʈR ���3iWȆ&��Ddw�h���>��fq	.�T6�e���2���t�c g�C2�5�AZ�PNm(\iQ*�@���\�y x���`A,��`�z~��"/�t���<勛�1bGT�I��,e���è�Y�J
=$�L�W?�S?�� jX�"(��	 �Z�cW��L�Q&`����4��vuSx8�m���2_?�<�时[@lb���i��!��8=�HF�^c���z
�.�$f�����q��Bw"i �ؽ5�2yQ�u�U)D�8�+"�0I�N��T0�g��.�f'�	,��i9D���ƽ}:�]>_:->�C��Q1��*���;��֔��&������"��2��
>0eHr4�y�0�4��&k��e[�y귖�0�4.0�^����m(�4��be|0��zٚY��O���*�;^���������?Jz��===#�٧���i)f@������3K�2��@|^gc��{��$S�v}cm���ť��T%��RiO8j8�|�����1{��\��ӈ��`��cb�\4�����b�>T5�ր9��U���g
�6�T�t���u~�N�����g!�,"W�*�=B� 5���Rw���SQ`�Bs"`0��8�ƅ:�N���/��+Qt�c�pݮ_�p��㜯R?VƟ�}L ����E&]�bY�y�u1ږ')W���f��\�*O6%C+�z��a8R�&>\@�����Lay��pl�p�@���1HA��Q���G�/�$��P|/Ϧ��`�1��MD��3���Ht�b24�N�'�3��ԴR�{4|�M�K<�k?���9ϊ6H}��ƿH^]�� ñH��3��w������s<�T�$�\c�	��x%����H�β��3ʳH��
���p��̩J*/����-j��z)u��--{� ��Ԟ���6 ��L�k�{�]���Q�)9,	�0��d���
�����e�q��9�fӓ����xsZ����ą��Ș����T�M����e��3�v/V�u����C����Vn@����jB�!ʆ|�����\ը��d��"bp��z!��
���I�ꋜ�<�����)�np&�r��%��+� ����cBNs��Sd�xohugKw5y�F�����i���	^�q𭚵�<�q�:8TIR�4��(}�"+�c���c�pse�H�m�J	���S�v���)&��ԾHQ��&�Q�LO�_�^\{����\6�Sqi*�p��|����#*�;�lN]_�;�3ъڭ�H�� �"1�S�<D�q����I�=�K��Xĕ@�6W('-a*���[4Q.W�RwhA�AQw]���( ������FVD|7����@bY9 �������`�|�g �Iz0:X�He�n�n��0vV��#.N����R/$7d�V�&���i5�e��m"q¿�\�<�DT��뛂�:��z��f`�D��ҘD���P!d0� ̮���F���0 b{w�DP���7�G�<V�=�יg��/��"���^��9��?����{s���ï��o����8���#��X]�|S��:�$��>'C�h���*�S�����~9���/:�h���4����|��tu�r���*o��5 h��=��-�����\�(���v� `�5m��;3��|�q^��/���a��n+O�|U�V�-��sX�L�ng�D�<d���Ll��J�Nbz"��i�ߢ-s�!�¤h��(�XK�Zp�cI9��Y�ݽq6.%3Ι$Ґ�c�'�q_$Ƥ.w�"l����h�F;?ay�/^�D$��h"�u:��|�O�o�S�K��K�cXXva0��2ȧ�嵩a����F~3��,���hg�3�;�|7��"%�D�t^�)ng��Q��mIJp�=�^��ϻpT7K�G	�k#O?�r�10�w��
(��&�YE�h�|K�=�D~� @I�p�X�]�@��Z�
a�t��W���)A�BE���Բ��Ҧ�w�%�,��F*p����?J��t��������U�sV�1H�@0Q���"�V��h3X��}g}�Kz!���5�
yLç���K���!�)S�/k���|��8n����Rw�ΘO"p�'�ը�n�����1m��7	�Q)��8�m��.ż��$�c�.��'	�R�=�$�i��H��m��3Ą��/�����SU�܀��σ$6����6���ؐKF�w�7EQ3����9ܞn�J��SC;߿�����f��c���|��~֔ޱ�8��`mD\A"�Z%rv0������Sԃn�U����Y�h0�7j�����l,3���}F�ǿ�
� ����o�9�>�y�|�c��e/[V��:��h��py4֐�26W�J��팄7�06[�s���Fh]�@X�B��N �J-�c��qw��9��x*RR�`�qG�Ϝ��T���Vc7.�y�a��!}�Ps�P
n[�"�"pd)�WFT�3. ����@ő$�R�ٜ�i0[x���,�b�p��P</�í��8�Q�,3��O��B�9"��U�2 ���⭺��j�<�W/�U?�+!Z��+�G*����٥l}�AN�P�4��Af��(V��ɮ�rƘ�EK\Pe6��|�&�-� ��H�����Q=F[W����2�X��Pt�:1�F(�}:��j(^i���@�>�� x�,s_4��j�2��Ytܘ6�4Yc�9z��Wʔr8%�yO��E�d���<���G�PR����
����"�ՠ �¢��U�j���H NJ~��E�ء\~K���jU�v����'�j�eY��-Q��nl68j��E��=ęAj��}��Xn�b��^tx5�:z�J-U����q��`�Vl'��nb���)#1�<r��N�Q�L.B�Q�f�-���� �}B5D���B���ZJ�ΜOT �*��k����Vx��PR~�RV�b���%�^��9.P����G�����&W�j�&��nd��м�q'>�Q�qd�N�e�
e��2���t�g�&\C-ؒ���P�+h(w��*y!�¤%y;`шqp�<*��a�9`O���"V^/�= ���< �5��w+I#�le����.��ԭ�
�CLӰ5?$���{�j��(�_p ����p����QYi�`J�%�/�bvБ�8�w竧s��������l��"�d'�!�V=K��y��L*��ͬ$�*�����l��BҶ �<��,�ڭs�P�)_�8+Xg�+	�NG���<�4���l��%��PD6��Ƹw��(-�bɤ^�ڢ����U��v�4�=ٝ�$P��9صZ��_���e#S���9t�/�&�F`�D��[�<��/�$ęQ"wަ�Y�я�\�9�|KwPzT针�D�T�\��`ǣ̞��'�㰿Q݈Z���e�w=�OL��r���`f;��Le����v3f#�IH}^BZ�'N ��lDvx�K�nȖ�`�fT@.+R�j8��:�I�w�[{����^��ѹ�`�M�bM�:�e� ���̉>OM��{*���=g���6}Lyt��,���N�l�U�֝":�,=�k*|fB��c�(�Uw r�SL�̢�M`�*x8��:=�-��}��fZC����k[��r"9p��㷵�?я}��L[�0�i�}&XԮYDh^u�"BZ'A+C\?"O�+?+�z��y8=BY8�5��ž�7a��*pk��W��H���l��!���
��$�|ʫ���Щ1;��M����N�����^4��'�{�fR37�9���4����;9
��H�DƺNb^�� ~"0�){	�x0�]{���NT3B[�W4=	:ȸ%��ȴcN̲s��ʎ�"l��J���E�*���h���*�J�<�u�,�h�Z 1ݜ��.�6gfB��k�����	*��MP�d��,���㖐�@|x�y'��I�+���Az�/n��=����`X��)��LWM�I��ͥ~�Qh8v*�=�Й�C�(��@cQn�b�"G�a�w��O�Z�cզd��fb��z�A-�E-O���	���<�O�����prdui%�*m�;�	�z�#Nn�(�ܛy�3�&�2�w��QF��k��"jܝ��^�}�f�	�U�=<�'�:��R�ݷ�cA-��v�c�q𲾫�p.��H�wJ�����g������ȳ&�������l~7O(o�\�\����&��6���i��x�O������*��&l�B}_���;�SE�5��H�� .i6"�:}���q/�#��̈́�6��rQ�X+��Q�'�Q��s�B4�)���c�MA���]Q��CX��Ze]�@D���7�����b��� �8��­���խBVLI�A�X%�{�iQunI�Y01��><��/�S��յj@�dP�|�=����5['�Ĉ&�:8s�7��k!x�#�d�:; ��;���_te����u7!CI0nzĮ�s�F(G���{3��׿����i�O�,<�g���^�U�m���p_�"7ײu��*Ā�pRnê�/�AХ&?�U^�S��]����؍=�QԆ95�6)ଣ�S0"ӯW�.~��=�������P�|�t*�r�����pih�q�J��ѕ�`5�+a�������W5���v����g^�-���<Ÿv��+5�����V���3�A�J��nbȊ��ݸ����L�1'J
�b�(����zt�s�&K�����X�Xf�Z��7>��.��x��6)�k���$�H=B�_�k.R��l1N��n�F6��y�)L�҉�$�̾"
":�0�|��o�f�K[����XGj0#��2C��߁ʹ����r�#\���h"���V�'7O�*|D76���V,�0Q=F!m1A�XZL�Qa���Tr�G��#J
rU�/0���軀
����#Y��hR;��8Q�~���@�u�sfXFޯa�ECLt���bi)��jE>A���q�!W�� ��,���#���zJڷ/�<��
���N��1>@�@�Pk��_V	)|��z������r}�j��Z�L^���	-O��R�J�s�9�r�!F�"���U��!	"�c�Ȉ踉�3�z-m�0�	kBL�t�h	�. ����? c�Dݿ� }�-�x,�$7��gK�qk����1�ϞV�Y$��.	sܻ�M�;ޫ���jk�f2͒�*�E,�g���P��]UnĊ?���2K;����^�Pf��H��8����~�ܱ�3�ء\\��Z��rQ�Ŵ9;��W�X�i9e�`o��hKCjrX�o����k�e��F��{�e�1��f�7K�o6�K>˄�|�ɥ� ]�Vը>�g��u|�4�2�=ZJ|M܌����ɩ[�ڪ7!h���@8�IB�8��)aX���[���l�����x�s��{��GL
��8Txݬ���.�a�@G}ׁ&���
�"�"���dM��W�-�3)���@���-SV�d�ʹ��ik�2x�w�'��ˬnP����9Q��o�^G,@ۼ�꜒��_9}�1UA�^�2��(c��!6<�
t/2p���Z���B l�)�*�!s��G�WAYKPH����TOf
Lt(yw��;��J��s�u���\�U���E��-����p�1�,���/��(��]'2������.����e}��O}E(�/ڦ�ک>Q� 3��szг��%�fh��� �4��߶4�K�Μ-�-���˒�TЪwF�&�7������
���ݰ�;&��i��U�Ϻ�L� �Um~�����\�K�Vb��U�va�)3!�`�9�Y�JݮA�lQ��j6���R���Wd�T[ē�F��	���xP˒z�e-0��R���r��Vg�.��I9��4�#L�7��(Ndb)��Z��f�T��޵8�D�Bx�Z%{����׏��k��U���x�edPmr+R�k��U�`�
�;�M.K֏�U�Ĉ������lW�,�&oըd�.M�>f->��Sq����������C2�W�tH�:g>�nC(q6����P�)�(���*��ݝ�yv�~�;<7HM���0`
l��=��/����<[HD�g�wI~�,ed$����g�O��
�6L*�?�tZ�/�j1�(u�z �&Y�3�`�}Q��4`娷�*q6v+�>8T�����?5�1֜�H�>�l�r��_qp!E�S=��̔ۖ�����e��$���Hi��g��B-k� o|%��c�(�u�+\�)�8ƤD�&�bN�g����O��\Ҏ��&N�N��D�MlƳ�o�3;����yה�Gr���"��\����~��UT���p;4�0�� 0e�����Ư�*H2&!����6�[�@��?;��9���"�w�e���N�a0|fE�zϝ��c�rԏ�B�q�h��ux�7l�z�|�u�Q����=ٻ��Z}蟦f6&L��F�a��3��{��o�^q�b@U�Z�7vs����>��T[�R_�j���u��[�{���ʹ����`���b�k���G�[�<��ܺ>J��6�ݘ�P&sRg��6Xd|t���̫S N�t�����r,X�5*�mzB���c�w�WBSGr�����`��y8�:�k���q������ \f�e��Xp=k�����?Ly���[L��Z�w�&S7Y�v�u�mr]+��B��\Y~�OlR�+��z?.r8ȡAt4��n0řMa�#tp����lU�H��𻇎���D��޹$<g|e����`�1��vMy>�iQ��>*:�˹4W�l'%���j�R��%�i�إ�����Z9EA�H�rtƵt�^eU 9�{�D#��󮢾8����T���R%�	��x%S��~�Ѳ�i��]�y�塌��*�B��#K/�E	S·�-u����s� ����6�̕���k	2��S����iUԟG�,?�O�����4�ƌ�s���� �Am�j�׮&F��D+�]q���`��y�M����S���v%y$��T_vC�R����n����]�����rC[�����3�d��rbfCPz�	����m�	��\ڪ�)����p7�r�x�%���vw��o�Ni�4�7��6i�ew+��Fa��#���8��^�T��wí�)<��@:.g�R��q��% �X��c�P-�j�p�X�H��xJ�r���o��xb�F��&�3������/��*�O����{\����9G6��i�܀�
��"&����*e��l�G�_9I�;��U���H;J I�["' S���qj��A��ͻX:��l�'#b��N�y4�D9�R7�^͜A�]�r�^����g�8��D��7"�����bw �g�����V�9��EI�r�X�٩�d�nn�À0���YjD���������|qd�j��t�6��5	�ģ4#µt�e�(��!��f�:�A�����zx�Ҏ3t�P��!~��0	5��@aF����ϳ{N��:�S�\���<�lI�ͩ��l��(�/��J��T���A@�e,����å&l%��`4 �a��	�]�L��Z,��4cij#��g<NSK���><~�!��xW5�r��Gɫ���A:�tE�|r�������̫���Qp���q�V����=��m3��5�>Jѱ;�಺�^����X��1�w+PE�r^�V�5��n����9,n]"-��v��cxlL���J��{b��3���,�f�s�K9�Z�G�L��X�{Zf'V�W��W,6$�@�O㗐�]"�_��.-�tll�Ğ5�F1�RyADz���$��"��:� �|O�Ro&��Kኚ�X�7�0>��2����k́�S�|���t��Nc�h�x6�q��7�n%�P�DrL�__	��Q��bm�7��s8b���2ѝ�T��G?��#E�ur��0X ���
Ѿ���mY��$h���3�~U�L@��^�����ފ� �E�t(O>��߁)��E������Ҝ�T��f*,��`����RJg!x���ϐ��Vk�)0�1yX@fp���(�Vd����<��1��A���E�;��0EL��%���R^�;��e2��#����������,��ʾ"&,}��\���Fr���4m���	?���4ɖc}y.{����c�zV�	��D�̳pS$����Ц��̉����c��ł�h�	�.��)�Ϲqޫ̣��V�%�֐�>�m�E��U�o��n���{Ȕ2W;���s[f����ٝ���E~̴u�CW��b#\w�tZ�@�r,���t�j��"��d�0һ9*���hf�j��4���� h�F����Р�gRo���>��+|P+ԛ��VЩ>����0��4��2,DJW#[��993�5[��ܪ�l_h���@ST�Bu�*��P��Ed���g����gx����r�G����&T=p��`�.��aI�L}�N��)�
d
>"��9d�m�W|'�3$:h�q�T@;!oH����͏�i��jx:s��"���&�	P�Է��s�ym�c��,{���l>�9��U�� �M��+����<޼/ͪ-�'�ZX"��D�����"cAA��dP�E���Yfe��(��{�8���h���N�5�t{\�f$��*oM\-nݼ��e��?�����#=&���L�2Gհ��)U�I�4�<�E}�!��|�(�i���>�� ���s��:�`B��A���+m4��L�/dc���w:��}n�;�ǪR ��a�;߆���?�
>8�Ș��V���n>U`T�� M}H~����|V�ȟK��m�`vv<K�d^����[����X��i�&ll��j��$��-���ҷ�X����<�s�r�yxk�z���-��ɍ���Vb���QE��I�2#g[hݳN?��¦0��f����c]���D1ͼB��Z W���b�`D�k���CnwxT��P��RL0�u��P���l�.F��ưuB���
���:Wx�&J�d(�ݼ�z�>ˁ�q���jI��[[�]2c4Vt�l�g�9C#�P�RqRP>G*(���*J��x��y�F���%n2�����`���X��/��;�\?�<��Ɣ��I��leX��dS�ʪI
�]�LI�^?Z5��ji��(0�) ڼ����;�QϑJ`�ԁ�%Fv�nB8�	��U�4��w�I�l3	�Z�@!�O1=�fR̯G��B��@k�$��jz�b�B�?� *�2���ڣ�Y��g)��[8a��!�N�f}a�jG���W׮�[��zDl%�Ʈ~$�n]�k.�����B�������7��s>8�07�:�+<ӰKu�{0�e�H�#�MJt�%��&|'���i[�"w��R��o�����`�
���E���G�|�3|zJO��>�P�ʅ��HB��l�����5u���u)�[��=�G��Xa�:�f1���H��H3��<�?��^����R�����vn�|�$���H�TvllRڦ�j��2�� ���{~8x�Qd�Gx`�a�bCI��zZ����3�>E>�֑`ј�wA�/g#&63��t3�L�F� N�b��Ǚ����,sG�*r�zB\i��@�wV]�SB+8�S�"`a��82x4:3*=�y���̝�4q<aCT�(	p��q��!�?ǂ�v�RL�9��R�&NR�Y��:ubg�x\8���Һ\�ݎO�?+�)z��J8�&%�P+�t��a*��p=\�]���IHr������m���$w�4| �
���1�2TM4��܄C�ڹ_�E4�ou'�j����R�~�������*��o;�9���HNe|ư��^nj$ �c+�_�l�nz���$�YTi���M6=	��%JѴ��߲i�[�D������j$۽ݨ*@����g�`���2?rur.��l g$՞�\6S��}bMk$����B��n�*���,�3c��ZC���������/�!����'��Ҁ�I0p��\m�����F��U\�B�`M}MM�C ���1�v �+#�RC�!�6^Ln�-�����S`��m_���ٰ�d��Fb��z��H����TЋ����U��Z�JpR&�rZ�w%�0@��e=а$�Ndf=撌$���/�(�w�d�F<�^������^	H�+�˱�<��:� �Ru�۔�)Ǉ�m�c�O��tHUp��Hװ�Jzw���o��'�{���&����Y��Kd��DO����\,�^�\�p6���i;���[�=��y0�*@��l�l�_�;}���k%H��\ d�)"����͢Fq��;�l(�(FpX���ˇ�'����)� 4������Y��Ab7�]�F3�y(��P�/�fD-5�7��0�~DbjW� P�m��Sf��~���a�I+ĲX[R��_I�n��G0�Z��t���%�iά7��؜d�Nr��5�5�5�
Bľmh�0����P4c8�o댈:�����Е��	�ƅ+Ew!�W0����-aF�?�a�b{iܔ׵�'�7,���^M<'�3��a�ǣ��?�EY����.����7�Qà�d����bE�:�+�I�%]f��N�@�&8�/���0��"�6Sf��M6~�dݼ���9Ö������}�t`Flr�~��ؐ��%��!���yi��}������΂�<
5��&�����M��^�k��9̸��+k�E���Vey���Q����nX�+�M0t�]�L�	J ��b�椤4h���w�s���µ����X�rxZ�q ��㩒�Q���m6��Ϊ�*���xt6_�&�.fl���9�F,pey�~�Hu�$"'�" ��:��"|���o��%K�ښ\qX�H�0Y��29���F*�@�d�W��宦���h��ی��7E�B���D������3IQ�Dmz^���6���0���T�-G��#@�r��0�{n0
�ݷ����Y��h���.�"~�Է@z,�������e���g�tø���|)R#�E������|��X,N���<�{p�JX�L���:�� D����1���@�=��[}V�-cd�B���i�Ù� D���s)L�G����T��������ت/�s���"�k��#��ӿ�p"�h�>P������p�HmoL0	z�0��5�^v.֖r�U?c����������ԋ$m�@����'�)�?�Y�}�Oͦ��к�1���T�6���G�ʸ�t���ju��i�E���G���
�*n�����ORg;0�&�Tn�f�A%�#W�M�u~�t����͑�\���Zw�Rr�ݴ�;�����_/��$���R�h���jhY/]����țj�F�i���ϠQ�Hm�6o,l	>��|B�$�6�V��:�-i���4'z)2�j�J2j�5�&�Z�[������[h<�`@n�B����߂���!�4J&b<y�J"�x[���G��\O�Tx�֬'�.ן)a��2}M;~ĭ*
�
"e��d�?�WAR3����s�@��cM��h�j"[iᒶx��m�������Pm�����e���>��,���� \��g93.U�{��h�������<Y�Y/hi�ՀZ����1�_�������A���P~5��&`f�\�(���S�m��'�)-��}�\!���',��-)M?���f	W��r�7>�?���Z2��)�����d��ʷr}�Ňśw(/P��n�>�� �
�s�h)�ۡM����IUM4*X2�*	��h7��GK��D����K�-��T�!���z��
��-�SFl�qj/�_d�U;�7��C. ���~��V��ҭ�KqA�۶fv�"����;7/�Vʏ�^�$l�pj-v��(v�J䴷�v&��j���^�-��x��[znG-�8
��xHب�<V]�Y�`ǰ"-#�k���jN䯌�6�S�2f���\����DL�Bn��Z�R~� Z���k�%.����x]P��GRǺ������?�q6.A�����>�;���W��&%YMdc)��t�>�I�qu���@�΀�<$2>1�t�&gt��Cw'��c�P���(�}\*��e�S<�y��ՈB0x-��r�>`�ݐ�s��/���7�<ф���x�
81I4B-eګ���/G�Eٶ
�[�L�|�?�����j��s(�| �rJO}�07Q
V` �� ϑv�8�TA���@+�V�R'G�	lο{�Uem!��=|[�����ʽ���j�$RY�~���]?gB�34 �[D�)2
�#ʍ��)0�L8��Ƕ	ENX� �������R�ˮu�0��j�DƩi��ɧ&���Qa�=3�����'3.����	��
�v��\ְfSܲ�k�e���^��A� *�&����uns[F���,v��� �J%�H(b�� Ѡ���}9|�ANz� ������*ǧ�S�����8���6��nI����=���ٓ�Y�գof,���]i���@�3�de��	^���؄���y�viWϩM�ő pT�;YRUY
j�ݏ��=�H�{y���o�Ԉ��`�"b�F�r'���89��[E>@�z���A\��g�k�6�rtn![���N�p��f���SD�,�ׂ*�tgB7l��ٞw��S=袮��`�	8M�~:���\'��6)��5\�^��,vp�h���7?B�Q=�L�ˤ:Nx&I��YU�Hu�^����֮\�\O��C+	�z� 8>�������K�O��ae�p�-+���"~�H-�����wr�r�$�q�|����`1LRM�n�ܟU��4���t�4��'[�݀�RD�h������-��J��9�whH�w\ƫ u^ɏS �4?�z����eL��+��_UT[��Hg�	KYy%ɥ���g���	,����OU�S�۸�U*����B�{e�­��uM�� xE��#~6x�|�8ԕk?d%�IɖI���Y,u�ή��&�Q�������{?������.��f��Y���T�����`y���ߚ�TMX���~D�"ƪv6�/Sn��d�Cԟ�Ln����Ӌ��_y�h	�`?�ՔNtd�)�b\�z��N��֧���w���f�`�"��pmfr���%k����s�K��N_�A��4��d~z�S�w!�F`�����n;^UW�w�����<#
�:$�;RP���N"��Ac|n[��F�p_� H�TJ��d��#͙b�h�|�d&�烾�6;����gO�][��\g����6�g�i�e���;�X�A��*�yl:�'_o�;xsJ�F�}H��� O�"�ըW5q�o׀�t��������X��ˢKV'��O�4=�k���!T��A�]��W��5��~wDh�Q7XZ|_�b�W� ����R�Le'���If5X��N�Z��nZ��0b���&���7·��U|d!RA�B��b5�,�����«M8��\|���Iފ���:L$|�lY�а�҄����!���0?�~��:�F9�{���0����`� ��<�յ��9��"{�͜&_R���'��;`��\��A�ÛL��'�֯��U���:]A���G��A��*  ^>��̓S��ү�~�ǁ��gDk���X��ar}��"t{!dr��q�����!e�B��}}�q=�H��ڐ��%5����'���Q�^�:n��o����+�S��h�OV@�1��0���nS6���	"��aZLإ�J{�b���oR>�K��s�������§�X���Z\�6�p�̸ͭIpG6%��"ސy��r_��.�f�l�����$�F'k4y�ؖ�i$=�q"{�+:� �|ż�o\^�KM����XDy�0t��2� �!���{�鐲4�vҦ�[hS�Iۧ�X7�{l���D�9������QNx�m5����T���Z���T#<UGu��#;rf�*0Σ9w�

��|UsY1(�h#7_�)��~@5sݳ��`x^t�@6���t^B��9')��Eo�J���Ғ>b�j�,�h���-�v��JY`����{Q1�߉01��8@�;���&V�6����{��7Z������aL/���3�h��p��+g��J�¤���ْ��!�Ӻ|"����c���<��hmJ
N	�vV��YŎ.1ʡ��TcG���LᎾ���)Yx$ؽ�Ƅ�ق&��� b|��Q�����l(m��>�@���Is��)f���e�c9�E�n2�iw�In��P\6�
�{;K�ψf����OȪ��+>~�T}�����Lؒ\���Z��r��1����(r6�Z���q.\�E�kh�
j�	�8O��XY�6��F����v./�����8o�gJ>\e||}���ѥ$V�3�x�i��_�4B]�2"��J/	�p��iS�[��6�Hc�h�w�@�ЗBk���CR�6ޑ�ϭ�]����x�c��īG��7�pT����݅.�A�a���}H �Q�
Z9B"@��d�1�W�z03�6�'��@�0�~���[��E��i�xp����
���P(��H�onl�E�,�Q��k��9�t�Ur)�`<�R�z	�<��J/�|��Z]sj��z�Υ��dA
�P�z�ܿbf�(Bd�n��^�h��f7��\��r��I%�O-�E�0!޺��+ҽ��2l�\�5����2��b�<�F��X�2:�}s� ��(�C���h>b�h do�s�d��V!���T�܄�!4�鏶%��Û�^7`��+L�1T[�4 ��`�߼�a�u?�
�6���栌<���y�U������ �,'~|h��ѝ؍��K0.ݧVzv�
���m�	J�Q��jx�ߓol�Gj�س�[CiąZ�%�K��[����ɠ��x�$�z�d�-�����b�CC�VXW��~����#��^@NN�T��8�����f��S�Ù�iI�Dg�B�QZ�n��;����!�k�w���px�;�P��RB��t�4�uȰ �.<���f�=��Fq�/oWn4L& ˷d��:��>�1Jq�re���
4�MQ��2N�t���ge�C*��v�P���(��*���.�y'���ZZ(b/�� V`;Əӎ�]/����<S(�8m��I��me��C��'0
�yoL�U�?����j��(��s I!�ĵ��QE:�`�����v<ˉ8��<�����[�-�����li�I�P�!V�=7p$����8(���p$�S��:�X��B>H� ��Y�D��ڙ�ƍ�Yo)k�Q8�Jm�I�N����'փ�+p���l�P%���z�D�4Ƥt��$��y��ʾs��Cu�qX�bN��#3���eEKء�=���+�q�e��H��W�/3��"&2���0:[5����ҥ�{;EąVv�{� Ie��q���H|�oHz@�����@�,�B�����J�����Ƈ��Q,\=j����υ�p�$f'�H��������3�h��5��^�u����+�vd$��ڹ7�L&T�*�R�+j���&����{tH���_e���`�5b9dnM����i˞>;��G�x��wbCguԦ6�kft����|��NОt���ݝ݄,��*h(@B���w��#S8���	��`���8h��:)}�7��R�H�j�EW����oupn��#?���,�QLG'��i�&DP8Y�auغ��7����r\
�KO=��+q�zP��8������!���*ZFa��ps�z�S�}BH�='����[�v�$�&�|6^���Ѐ1��oM�Ieܺ��گ*��O��4�"'��Q�;�R���#_��)�� %�89�BGH��Ʀ�3^$�� j%����p�dq��ɦ���+5T���C�-	�ɹ%�!��Z�_`���N1���[�۳�*����T����C]�(bu(�@T�M ����
56ӿ��e�kZ-����@�$}E�P�~,ђ�Ϟfᬁ�e����/���&��U<��@��,��6�U�����t�8��M3�����zVv~����Ѕ��C'�.�,��n�ج�b��c������OAd�Gb�,�zh!��1�¯PI�����ڻo���'p��CrPC6%F���'�A���ZNZ�B�H�ϨRI��Hw��SF�ݬ��G��	�U^�Ȃ���AO�<>@u:��R+���O�1�)�8cw�L�*e�p�=H�.Jp���`����*��O&��վ�΀�-����O�Ge�*\�P���+6�<i�ٙ�;;�s�8o��*��
lu�_
v;s/����Hl�Q �1�"��Ճ,Tq�ЀP����!��޺�Xk�h˽V'�S����4xV��#(O�A�]=h��x��F:���LD�!b7�^{w`�b x� �'�.zG��k����I���X����U�n�E�0�������m0�b#V�d�uH���G�5Gn���?��&�ڣ���H��l]�,:��,�'&O��Dn������Җ!/Rh0ڠW��g�F����v�{�ZQ׫�s����;��<]:о�1Q�}rLY�ќA��m�h8�%����xÖ�6�Б\�p)�?�]t����+|��%�{����4S����C�~�J��)F�eL���Rɼ�}�re2t�dr�Zq�q��\N3��"r�������F�����{��om5_i��b�����p^�)�i�Ӹb/�+�$����Va;�01춍�nN�<������L�a}J�K�bd$W��\����5s�z��k�`�}WXҠZ�f��J���[��,�6uh�`q��4IY�xW_��=.���l��oL�F"��yRS����&$X�"��q:_0�| �Fo���K3���X��v0�c�2/�P���5����M2"�'�_tqh���6$7;2�i��D#{�091�
�Q�s�m���Ē�����b��T^�1G�7#6b"r��S0��ST� 
�V��W1.Yl�h�u@�$��~fW.@��r������[���1At�����)�E*���9���!��l�Y,��1���q��Jx�yR:� ���~��f�1*a@7��!�Vu�Jڬ�QE粔��3��FZ�L�����A�o�jl5����ݪ%%�,2h��Yw�ӵ��"7E�ഗ���]�f��m%��	�p�W�T��.�q��zc1ݲ�z���~��d�$�s��#M�ݤ���c��;�ÂE�ɚ�Cܧ�ϊ���������V���"���(�E�MV�#�@��n��~�0����;f3�J��fd5B�������~�T�T�*�À\�,~Zmq�r����%���I��U����XU� �h�7j^ڈ/y��4����AF�u�у�ǩ8��"o"�w>7�L|��t�lSCV�l'���a�"4]`e2��J�d8����li[����5h��`@���B�>���$[�qڶ�j1wX
� �x�:����G~�G�T�� �]�u.��aZ��}�tf�
Հ�"��d9D�WMԆ3�X���M@l��Odv�g� �:iW��xa��.��7J�P�<~�4��Kn���,,�@�V���_9��*U-�����E��UAN<��/�h��bZiʙ.�\�/�������AEEkP�����xafv��(�G���P��ل���(�r�E\WX>������-�
�Kgֺ\�,Ҙ�m�\�������2X \���eȚ�Vʭ��}NmU;:�(e�&����>�0� ��s�?���&����ܿ	�4`�e� ��� �Gy� 3���>���m����W���p�
O���[���.k�U�JU�u�8$! �*~w�
���H�PKKA�їYv͚q��.q�<�L6V���ݚD*l��Wj�݂6~����շ�i��l��M���I�x��Dz{Y-��]�>���*VS3��b�հz�#���١]N����sK]�Af�0ݙtIX�$�XD�QBd��Z����v���1��k��v�T"9x��PقR��Oʴ�L7E��)�.7
����������,��W�v~&�\2d٣��x6>�9q+z;���OB��7�2�t4��g�D�C��c�Po`L(��*}s��	�hyb�}�x�# 3�(^�`���ө�!/�O��*<GA���) ��I�2.eP���#&G�;��
_��L�Ns?+7��?�jz>�(a� +? EС���Q�>�`Q1���v���8@���.�b!��/.��}l�o�K��!�=�c� L�ʳw����9$�m��/O�SI,B�|� [�s�_�%�8O��C)��j82����N%��r%��ͨ�H���+���:��D=l�Ɵ������O��KN�3t��LT
�����D�t������\���#c��BAej�>��
=O���&�h��%[P�L�x��V������~�������V}U�MK�|ҽjz�#L���
�{:��ݒ��	��P�f����a�̈=E�Y�	7��!2f"���8�M:�3�M�^�ǜNI2��̵v_�5F��0�T�9�RK�jZAz�a<�~-�{o �%�x�b`.��b���(ᲱG)�[�>6gE֢�,��G;�Gyg�\�6��t�'t�~3N������ɕx,�Wp*��B��ބO�2w'._S3<�d�`�=�8�I,:�%/��艍h���nR�Ȯ9�p)�(�>�?8_hOYL���p��&?��Y�u�[ɯ��T��>\E�hO�,U+���z�S8�t(�dq���I�aی"p1Y�u���&cH��A��jL����Q��$(��|������<1�MeDe�����*���*
4C��'�����R��	����D�i��� ��91.zH��ơL�^:� %6�����ߜ���A_��!�T:�/�>)�	Zz%?����m9������FI2��Q�|ۮ1*Qpo�&���A£#Hu�!��L 8Ξ�(6.�d��sku��?���ԋ�w,�Ϯ��p��%� ό���0���a�V�����ӗ�Nw�I��&3��C�MÜ��G,�XO�v�m�e�@�~CB;1���Onb�-�I�k$�!�^OӹD�
�Qd,4tbRe�zCiK�l=2���N�~�$�-���{�p�FUr��w%!�E�b��ЁNUa?��e��E�
�wp2F�{e���ܤ�^�\ʑ-���B<Y��:>R
:������hcrz����pտ>H(QJ�D��;�j��u���9�&���j�A�|�����O���@7�\��I�-��6�1�iLn���Z��·�9*��l���_�;�;nӯ��I�H'5 �3�"Vc�^!�qVp��냱���k�9�X&�	��'����nw4���JeqAss]�(���PW����'hD���7�̔r�%b{�� �s��I=D�B�E����I�w`X,|T�P�mn�]0�~���b���U�=����WdW���������5�����¡���~�|���}��:��������4�z�G���!j$�0u�����IF鷺��{��{�&$�ȱU�v��<�����IT�؉����\�<��
e�a�@�Q��w��Ñ��Mz�L�M��n=���d]�k������"� [�-�S�IS��Z��L�~[��dD�*��}*�����-	�t�7lry�|�LbR̗W�xS������'�����8Ǝ�9�5:b�ѝ̀�i^�8��Ĥ���e+���^��V��ZO?�Q�cnI�O�^�O��L>�Jq�Hb?s��� ��ls����"�8'"X�g�ZRH�D�C���	�6�λऐ�*�_�`.��ZlXO6�
�:F�y��y�($s�&"q�::�A|;3�o��&K�8�maX�:t0��52�m�ת��(P��O:����dhɧm�ݩ�7��D(JD^����n���Q��m������J�x�2=!�T���G���#1�~r�<0D�eo�T

�k�2-�Y���hY�y�>~��9@����*Sn����c�l�`t������)c�4E�Ǿ�T�|҈#��G��,�b6����lh�J�~����;�N�q̧��cv1e�9@�.^����VФ����F_�--?���	���Le��ȟ�ʡ�'�W���<���_�Z�m"���9Ӱ�n"��)�o��������m �9	+�mS��O�.����YlcL�̿�V�t'�̟�m$>O`�����8C5�p�ԄV�S���M�ul?�⦦�%�P��3Y�X�d���~�Y8�EsLj��������n�,r%�Ȁq�;����� f?���r��%�~�t���y��͒\��Z��r�Mj�`�-�^A��P���'������h҄�j����.���/s�l2�F�+�,����F�#�o���>��|���!ZV���.���74x�2��Jú���h��U[�[���hm��@���Ba��p%������sS!x�[��x����yG}�����T)���ڽ.���a��$}~����
P��"�KdtvQW�MU3.�����@'�I�������i��x�EU�������P���O��eI��~�,gd�����u9D�	U��3乊�⏍��0�<
k)/9�+|��Zė6�;��5�Q���HA��UPO���Q\f�� (�K����u�Tc&ƺ���Y\\��!������-Z�>�f����%Z�s:��4z�ҕ��GG2�N��Hȵ@��(�})qtv��( ����]>�O ژ�s�f�L�5��������4�l�����y���v��ZJ�'I���B�Mk��ݗ�k��
���ȄH��@����U̧\�s�� �[�~r~;g���Kfm�L8v�J��PKD�G��� .��UIl��Pj��ٟ����[�~��G�d �^��xת�z���-w�_�y\T�y��VN/��rͰ5v�#�EyT#�N������$g�f{�����ֵ��D��Bߐ�Zl��ُ�~�k{{����9x@P�R8��*�$����BS^.2g���9�o6��G�Wd�<&��d��E5>�aPq��1�q�\j��G�2��to�gED�C����vP*��(*�k����y��ψ����ۤ`�������/|���J�<�OZ�n���r+IE�negA�>QS�$G
:fL5h�?�w���Jj��(�M FUG�������Q�b�`������v��8�Q��I�_�J���o���l����F�!5i=����8K�.�;�&�$��O���N�HB��M ���zW�ڏ�c�rM�)��8���)+Ni��Mݘ�֏��í��o��u�$D���ƚ�P��FCWE�� ��ę�'�����߈����V��8�����g�SeE��`2�jc�mZ&�h��1�[ko���)�1�>��������Bѱ�g��S|�+�z6U䒪U�Զ�M�x�٣���I�Y�!<��Z�G= ���D�Z規�f0�n����3�P�+b^dÉ���K�a�vZ������g�T�hPR�0�j5����u�r{j�&ʀ��3jN`I
Vb/����:��
z>1
E��� �r���LwgkX6��=t�~̲��N�Z��w����n�,�G�*^�B�4���y�w³�S.Oࢿ=�`M�@8�$�:d����n��1D��s�M�'��VTp��X�YzH?��N�L����l&:�eYf��uN��`V�(�c�k\��YOs�a+���z-m8oy�� f̟��Wnaw0p�b$�pc:�3+�H^=`��<W��,@$c��|lw����1]0M _���K�ڥum��V4~��',ɋ��RUTc��W�_7���c�ۺ�9l9H�oƜE^ڿ! �fӓ�K�Z赾�W�8�TՓB�9�	\
�%�x��g�Um�ʰq��S����t۩�*�K���l���_��=uޱ��  �2��8W6��x�i�k��Ǻ4��Ԡ��E,F�"��b��b���s��"�ފ�G�cw��׵�ɳ����J��)�A��.wM��,�/����Cvvn�@���\�C]ܟ"�Sn=a���4��
�Y�ǹq�����dG�hbͽz�A�������~�y�M�q
�F�p��NrFj�%��'��^�;�NPJ8���{��Ys2��w�^F�9��J��?�^�.��8ŭ�lc<t�:�FR�rd��zl�_��cm���:p��HCu�Jfɣ���)�M�.&�e���r��7w��gAO
le��\e���a�6�F-i�"�������e�'*��]l�A�_@�D;i�̊W)HH��� �U�"����96"q� `��;I��W����X�M����'��g��.?4�Y��E�A�L}]�	��H��<���D��7)Z�m�hb�f <߲�d I����d��IImX�t��K��nk<�0�uƣ�0j�p��{z̉Sd����f\�N�5�Q�*�N����Y@5O�V�
�xP_:]h.����mc���J���v!�J0�q��!:FJ��M�H{�X.ס��s�䱓�<�c;����3�8�
H�wm.�ȅ�<"y����Ì��쯃�Y����(�5��]҃0�:!8aQ!�)�1����S�"��9�V~6���b�<��x���r;�����t�r|r�w��'�]�Ҁ������Ibꂇ��y#+�S�ɂ}"�5{z�� ��$�^�g��۸���+�&��$5V�Ⱦ���!�캍nDľ��Ul�
0�L):�J�*Jb�ɤ ���Ns��%�!�ǀ�BXO�Z��"`^S�~M��e6u��p���@��_��/.tUl�� ĥ�pF
y�"�4�n$�[-"�xb:��|v��o-v,K�^���F�Xu��0œ�2%�u���,�1���J��%�uh��E��<�71�1�VD�]��fj��b�Q_�mf9���n)�����:TԀGF��#,Prw^�0��;�R�
�O��IY⍔h�R�]�~Z%@fIJ�h�o��*E�0tt/�4��0B)�T]E���o��F�"`t,:zg ��gP�J.f���V#���9�p�a1���@m�g�V+�2PH�:[A��c�������L 2����%ߎ��a��˃����5�������ӫ�"���*_=�+�#�\m�	f����ؖJ��.B$��AXncgi�p�ҎO��ڥv$ٺ�����ٓd�+WۄqE+�;��P�����b	���,�������[���gENkn�3�2�vwn��a9P�;�;�Aȗ@��f��� x���'~����
T��}��\��Zc��rs�N������X��K�/҂�vi�h��:jT��NC�	K���F��އ���=��{�o�>�e>|.ϔԢiV����nk��b�4���2�D�J�0G�!�:�Y[�ǐ�YŎh(�@��NB���KF}��2����NXE���*xG����LG���Ⱦ�TdC���	^.��a�}9.�0��
�os"��d��W��3��8e�@�
��ls����Zi�G�xAJ}�	>���X�PY"��jvp�fv�K(,�l���Zc�WH9�[(U��*��On�
���;<E�/ԯ�wʹZ�3��-���"����i�bA�!�P�a��JSf,��(soP��f3��a�ƕ�h��\����vJ6^n-H1��S?�Ro��N�[��K-�����2���m
��б+ʣ�}�c�X�(�w]���>sC� �]us���_���a��5>W4�^y���Ԉ��Ʒ�6����sӪ�A|� ~ߍ:�f��
���?�.��rG�Kz�U��s�� T#Z~m9(��iؾ�K�%a���|v�����A��B"��{s��l��1j�����S��6}Ƿ�,�������!x�Nz��-R�ɴ=+��wVIK�e��|�#�#e�� N�g���U��/fvޤ�*�����D�zBZ}5ZG���v��g]�kv-0�
�x�1P�aR�������ݜc.-�`�w÷�*�)�b�:W�[�&��WdO�ݼ���>���q��G�,(<�6�²�2�dt��mg�c�C
ےm P廷(4��*s��ݿyضu����Ξ�x�`l@���Vb/�U���<�}!�	���wI��/e�:�Y�g�1��
��Lp�e?a����j0�(�V1 a��;�ᵂ�Q��D`����vMƕ8�;ȫd��K3־��3:Bl:���A͸!g~�=hn��6DAʩv�⇥�$>��R��I��BOE њ�ؕNa�
��Mws)��8h��ZN�C�h0��q�>�W��C7�k�Ds;ƕU��5�[��[�)5^�4_�`��zk�����v�	��̰�s���Re �zJ��Q�o�n�&C�8�a]�[��n�}�]�6��JX��L����ØO|�'z���������Rl��ˣ�:�c��}P����¡f=���e�AUf����.�ón3#5���W^?�<�čY����vUK��1�}�`T��]RAc�j%���rß��{e�����׈�L^`dDbb�|$�������:��>,� �X�T�-h�q=g���6z�!tZ���M��N����	�?g�,�W�*�SB����Ww]Y�S)����z`%[8��:�·���� �;�H�����3p��,�t`�?.�a��xL����|-&5�VY�lu	(h�1Ry">&�\��O��+�>�za&�8*������Ż��aQ�2pD�g�k�熎OH킻)��~�_�A$��|4���`�1��Mۙ����� K����4�Э'��<�,�R���TP 30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�/ڜ4�{^�{]�$Ht�E/Z}1TWZ�i�ˀ���9��Z6$�x���<�������5~��ߣ�L�8�6Z�^��3�B��˞� �Z�>~� Bc�wz�荏�`�ر1�y������P��v���cz���Q�ا���@�j�{��T�,2)��2{#��X�jEǁwNրv�t-+ ���2���)D���?&Ìw��K �ڀ�-���9E���YW�%����e�1�8�3��c��<G��Y>i���9+��=��in3�4�S�@���`�����j�@��I�`�39�Ǹbн�>D,:t��N��@wReb�T�
�1�掚l�A{��K��ү�!��'���^g}h�2�+����1�V"5K�AO���9�����sǑ9MܐxZ:"��?�_�=�h���G�9��eХVN�Ѩ��vdv&r���C|�4��|�C��>��0�� UpM9��!)!1Ê�y�kh���9�qȤ���%r����XX���|�(�LA���0;DZ���F�F(ן�\ܝ��)��h������ri��H �hf[v�Y�U�h�>p���Z����.����;��Jꋍ�	�!aH>l�#��wP7�:o�G��^�9��a��=�[K���N��T�e)��80��f�<�<��*0쉛���G��(��e\��*��c7ͨ�6ږ�?\���� V�AW�l@²��ހL��rmbm�?ɐ�D������P[X��9�K�L�ݢ���������(,��{׌�#0M`^�[���j~���b��G��_� �W�*��JPסs� ���-�gdxiN�E�AD�TB�~c;d� �b�%y�����_�Zx�;Y֤͙k�ֈƟ�]��ތ���(���Zcϋ���leY�yZ�����n'�b����uF�kS�8Q����eBy����Y�nFh%׎=���o���Bڨƕ�S���Z��[��!\��h�!��'�j �?,��h��	���[�������?El�p]5D��v�Ohu�4�%���2�Y���>�g���n5G.q�0T�� @��/cI��%~�~[n'Z(2��Y=s�m^eK=�Tl)�?aoX���:��0�z�0<�_9M�E��Y1K��0'v�u���Z���.�Zͻ	�>:�k���S��<�v�Po[h�Q���O�&B��6�"q��zF�H�r��7��G��yfޏ��Ф[��A-�b�����K�*��
�h�dݬb��@o��#n�Yw�����g�*
��R�< d#�m��d쒥���w�?|�a�����Q��˦�F��)=\�����`�=)M?ܭ�Q}�{�*M�#���c9+;0,[�?�ټj�����~��$=8�ܷٗ׻+�Ab�4Ԣ}&��<\z��F�̔8D�Y]�E���%)�7��s����Ō�5��J.�����sk`�H��V���*�uHC�����R�4
�����1�-p�GF�{l�z�X���1�^�g~�-!]���F	J)��Z��a���G�
��"��0X�A�fF�g+95@X�wk.#�"_A��K�Mn�����[N�d��m4�Z�����S��ʑs2�����x�t�z�m�?2��(?Be>���G3F��~i��p�_�{$[z�"t2T�Wu RCG(	�L4��
ز��!I��O��Te�*�}y��Eo���ͮDx^��5!xf����.\r,�W���)���b������<�W �ߵ����0��^lh�AUnM�#��qYչ�]ק �a-7�|�x����nblC�0B�\ó���$��1|�D;x��U0�ibL0�۸*t��G%%���7�<M>��k3�*G��R�@����J:ؼ��a7��N�-ϳ��S�w�.�����Q��[�A��8S�c���d^O'D�<��W�(ew�Gp8p�l�%`�c�ۋ����Hy�t�v�=�u�~y��p�z�D���a�]���4x��+�=:��|��3�	xef���Fʗ�O/�8�uj {���$�f�E�@+���iikn�����3����[C$DE���J���J��~}.�]{�2^6��%�vڛB���˘�̔�f~GTcc::Ɛ�S��x>�+��y�Tb��\�PT�4�,�WB�ac����!i��_��j�\HɎ��2� ��q��&[jT�w�
�v=8 'f� ���2S�.��%D���yMh��"H��T��g-�ѳ C��YQ�_k��[N~1�v@2w��1:斓VGVc1Y8E��FI�+v����{b3�4;5��S%�(���Q�5`s@���]�o33�������L�D��5�NP2@�ȧeD���1����	B{���E�+�鳕�W����X�hX欚~(u�T��Pf+K���Ĥ��E��'쭗9ǳLxY��IO���@�⬈�D���3�1e
�N�7򯾆A��՝i�P��4�l-��2��Q��N�P	3k�+`-j?�"�j�JI����� �Ё�Z
��*9u/�4� wϨ0���H�:�@`��,���y�`�ur��:�:�G��{F��hO�GW�&�H��g] �f2���S�\��}���OwŀTdё�J$���L)���Ca\� P)yH��ͨ-L������)��n�����z�q�Uќ�X?���U�+����F繥�2�9�VFrF��	�U��s�\d���c����5�w���/Bf�j�TKMI���n��D�>ћ�z͋���8eaXj%����|�p����8������p/Ƽ�z�	>��He��I&R^���A��i}�@V��5�*�٧������rg��,Nc���*�k�)l�d��\vB08hWO�C�xi��{�k�������AN3|��E
mF�5kx�H՝��v
��i�@�P�0�M�SE�
�>�F>	oۦ�oX��nҠ�q7�H������c7,J�M��m�zV$!3q����5Fx�&3W���E,	0�A�)��� �5���$��痕[����>p*�ӆ2J�5��W��4����wk��j��7���h�O?��1�ǎX6`%]'�gt��'D�wx����+n-�r���>f:T�����+�r�����~ӌ�~ML2Z�:�՟fpLFOC�u#�n�Z�#L���GP�'�Q�t&Kv�%at�"�Ia�`��9vn&���$C
���(O��Ja�5ӦRO23`B��4;�`<���Y� ��ɕH(uC�w�;��4��BǍ��uL`����V*��H��vmZhJ��]9宆�Ǳ2��G����ڍ`�礘�槁/����p�չ�� ����S��T�=>��b��5���R�A����&8q�1cn�M&C�gӡ�8�ʰm���V�ɷX�Ɉu���	�� \�y�و�QY�V��b;���h�Cև����{Q�c��Kz(#������<}Y��L���y�նtB����e�
�KX��j}�R�B��O��CN�Y2W��Sؾ��
�_yo��a<���d}`����W��\���kP��F2�1_�q�'*�d?�	/t�k���PY����a;�1�VvgO�b"�X���^L��"�}i�Ѝ��﭅X�a?�l�3�ݐ�8�]Ow~�5��� &�l
��=���F-	��Dr���S�?M岬 ��.���ȶ��W��$@-�r���׿"����#M���,��*����(��/@�QP�W��xmZr�$���q���^}O�=��&����~��#��ޙRok1���&�s�%Jt.6�&s��2�8���W�(��h�!��9s����2Y�*�E���qMU����D�,��M<,�qx�����M��LM�_���.�@��4�'�����ڙݱ?����;�i��4L!U�L'y	�,��Ty"p���H�
���,(�4ޤZ٧����xa�=m�-;�����-eF<-� �.R�3��������yۋs�����ú�R��壁��}��O��`N��-v\�졿C�ڑ�Sz���;�l�zI
y��'B�I�#��\��%zW�����d�Ywt�ň�Z�B�@��`�^T�f��aޜ��v�1@\��������%L� H�i�t�*Wb �U$8A5.�\����WX�i~ҽ�Np;��F��S�C��.D�P�L���g�&�S'M�:P-�m�,C&��<E̕1T�M�P-3^64�P2�u��Q��IRA�\�����~�R�!b�i�]�V��x7a�@��Y���[���ߎ%8s����}o�I���(��t�F��C*=9���]�Q��u�~�^t�K��-��Sau���O)"�'8�)C�A�^�$0C�-p㭕��>���;�Y^��B8�0��\�\w��b7���I8ƈ�I����"�J�6���}��9��H�gJ\xZWA�oV���_X�	�FK<o�w���$LR{�6p[lJ���z��_�;d�#��|��x }9�U���l�l��c%S��"���v.�?z�'K9�y�~�	"�h)��N��O,(���CE���J���o���� ،�r60�{b�iU�e�(�$k��
�/.K.2 �n�E�	��m��z/��[4{�E+��88Ͼ�,�ɰ�H�&#z�z�ߙ,�1�F+ɀ��)���F"��>�����АX9���Ibv}��[�y�k�fdEW�v.{�����N���%�ks>��riU{��|~��.g�?P�4@�}�_���)�)��Z{��� ����O�㜾U�_h�}�|�I�=�}����Zyؗ"�"�K�a:�U��]!'�[�&��/�K�����S�G� �c��˨<y�E]�T/\�4:Ł��2�i��	�l�`�<�8&������`�5e�&2����A	tƧN���]W}Z��-7�D?%����{P���kfǖ���ж��B��v�hVc�5�Z��X/������8A�ZŸ�����nJ J���+2�߽����x�w�������7yr��JΙ毚0�\Lj��=��8��/�'�A�N�w��Ƒ(
�q��M2��
�:�I���67� ����A2X_d�fq	;m�:�C�Fr���0K�>&L{q������t�93 /�n�X"m �OnKh��t���jN�\$�b%��f2ՂX��}�����Iu���Yaߓr��%ގ|�����������`*����K���ā��c �0h�-LS ��36N�Qj�\��r٧ɜ��[>RC5��
֞ȃ]}Bуf���\v`����7��[�*�X�(�D�!�fq��K��x&t��[Ͱ�	��a$ݼ����8o��u/�������δ�C�g���b3�R� ��]��AQ�"ҁ����R��_v��^�)�g������["�,'���r�Jt�~��__g�vl�oI�}�=��ldA5&��I�t���q�ʸ��p��Ț-/�P�A��>�N\6C�D���8��T�u��i&��ι�esi(an�h/7��H�dSm�
�,%1��|96�Yq(��M����/���e�P��cCF��ȅ8��Aǝ?;Ƽϐ%P�4�P=��cDϔ<�}35���@��ԟ�ύ��J��!��`����2\�jj?��УE��z�n;�M�}64C��|�iQ(��*{;vL�Q�kzI��$�6�3���HQ�g� 	�(C�1���px��̬m���]����	O�V��+�P"��4�(/J�s:f���5]f"5a�/5��.AI�7��v���Q�[y�O���c�g��D��eA��7��=<q@��t������.҄��D8��C����2�������7S���V���㊻�bMw�4Q-��ߞk��⌺��O�����_���A��=}pNL=x����_������;]�u.08Z.��ǿ��.R��3�P��s���ۗ<r�5���#{� z<�R�Bʷ��
d�y0
����L<�:Ο�������W�0�֔y}�:�ȬZQ��>n@U�"s[��g��iy��ž�oKJ�1��C�Sn�:Tt��n�낟 <��7%R�`��ֺ�S���؜����Jdn�-v�]n� `;d�����5)Q%�ź
�S�D'�-�!��J��+i��vpi��ϟ��9��d���k���f5j�1�ؗO�Y+W������V��	��W���<�1�/{-���Rn��ƌyṜ�&����yֺ2z���м��nBx�S��|�Y�ޟ�U+�:li����@��@[��$��f|�{/���{[�m��j�Z���\�"~�%	0�ޤ\Z���g�z�fn��ov��&B"���J4�!TӞ4N|���&"Qoޠt����n� �6�I�2(
t�6|f>!�aG:����A+�7_��I_s�K<��[��CO#1�$8��U�=�������*� 0���N��#B?$����u<�4ϓ���3�>��0tdU�O��v�!�
��a�Nku�(�;�f¾�:���Xβ���G�X%4��/�����7�,;�OA��gAS�v�̤z�j��)"/�h�����rN[��5<����vE�U��x>�f�gO1�t���U�(���@���zЌ�.�>ك#\BP�To�3J���f93�I���(�b݅�{���aeցh����S�Ͻ�H�*]���hh�򴛙�5o�e	ͮ*9ˀ7�X`6gD�?�����E��$o�Wưa��]����L�&�m�W�?�̃D����Eu�]ċSv�ژ�1L�ǐ�y�����j�����I��^@�Z�G�j��X��̪���/�d� �Q���M� 2ꡇ�8�7~x6�=Ea������+�1�;q �#�%�@�&�%�^SZx�;f3�Fc�#]���'P���ʧ:r (rZ�[%��2�l���+����������ڬ�%2���<8^lR�`vBSGB�Ԩ�Yn �F�T�%��dV�o�O���j��J�S�Ͱ��T@[!\�xL0�4� /5�?y�h��O	L�P[�ݓ�����l�~�5�ykv��hb+q����_�3Yű«��v5�Zr�}��? t�\;��F��땻'g�&ԧ��s-�R�=x�7��^�Q/aܯߠ�K�ݟ��}��L�����������K
vO�)� �o�T,�.�+���S:4�@��X,ıԿv��[u��|���s�8�#-.q�.�çu�H��Th����Õ�&d$��E�Бx���b	��ݎ*O�@�_�8�bH��o��n$Q�w훎�~vj*w��_�t<��ۺë́QCP�d
awέ|d�_�O�#��Q˚Q��3�)��B�^�P��ުK�?��Q*R��w��#Ʃ��+@��,(���F���%�*�9MM��l8�
��$�e+ٞI��u}���<idH�+F/n�81��][n}�"`�)�8��b{�s�D��Nʂ��7�4֘1=�`�E�rr���n�"��C�um��W���E���&�z��13Ώp�h��(��z"� 슌j��z�~��	]O��Fv��!���o��i�S�@�
i���a��F��+F�+Xg�kw��a��oA9x�z��Ѕ~�.f�q 8m�4��-ݠ@c��W(s2�Y���c�����ۇ��m�>T2-o�?/{(>}��G`�:�KT���TJ_�M�(��o�T���u�b�GU+�L�噆yjؿ~/!�|��x�TR���ʀ��D`Ž�ޮ����)!%ڣf�{��r�f��"d��dE��i������K�������������%Ā4AM:�-�7_�f[$%��@�-ĵ���������b��{C���	�!�GO������|*�A=P0ZB`b�����t]<rr�/��P����+��д���Jb�@�|�3��J��?���[a�=�N��-��Y]�`w��x�J|�Ξb�[�����K�c��Ld+����q��Ω(ЩG��Yp��d��c�_輁P���&tҪx=\+d~���p��[������aU���<�䫸�=�*3��n�s�'^�@��د)�"�/����"ڥ{���$�u�Ev�X^6Yi}(F������x�Ὑ$1���Xt���%ȕ�B~xWo�j�b�߇�6��+�c#nBBd�����a��~�K�cG��.f��ԡ���y���q�P�����*����D���9E�����j�N��[ �22#�Б�4g�j̪�w�*8v�U�T5� �<�2�L��A�DX���Ơ����ڭ�8?�Q�4_�� l��ėY�~f��>�H�A1]o_ ���l��Gc��Y�U���+c���.P�3?|�4a:�'���'{��|���5@ !����3`�̸i{_��D��,�G�N[�@���e��"�1;1Ҩ�S�={�p����6�4�l%��n�T煻�h%����$��aY��1CKF�}/�|��wg�z�N94��x!H���r�� q�ϴ��ѫφ`L�e׬jN�m��ˊl�Z[)�#M������%�(Ǳ�	�N�3x�l`����Ǘ�W�fI/'K�1�� hgD��z��+��u��g�M�j����խY:�U��@}~��ɛsu�:m\G�5�F��,O's���4��JCgj��,
�ۂ�\�L}��O�͞T1�p���R�7&)�?�ꐍ3\Ƕ�����ѩ��u���j�;D���aOĘ�&u�'b�+P���{CQ"���d�f��T�����<^K��P� �u�w��'AJ����:|�e�0���6�`�n�9�G��Kd�x�J��uq.c��K��[)�2�x^%s�5��L�H�I�p���^��dU�_
򶁩5�F_�u�^��p�����Ȓ/�H��)"��Ы'ì�g0^��hCto|pX�Џ��V���	Y�SB�7A�00Ÿ�����7���j��Ɲ��o:O�i�.J�ѩ��~�*�垃���"Jq�yW��tV'�_M�����qS�w��$�6�K�nl��!��p\_�d)�α�h�M��9G���&glI_wz�[�{��}���t(('�59�~�}D)�+&�������xX����H؅}'��� �}�ǒ{�b��>e-��$@�1�);.`�� ��Ef�B��yYG�zd��[ַ>�)A��^����zǾ��Hzvqzܼ��n�;���x+ޒ��������38`̯�_8X���Mb����Vy.�*fY�LE�gS.�����^p�è��:�s����^V{^�|{.�T�%E�@#�_��P�X-D)L5�{�UD =p��8�{��9eU�▒�=���#�����{]ym���W���6��U(��6|�'U)�&`(c/�Z���r���G�ǵ���4��XG<.�]�]$/���4��E�ȧ��>ut	RC��u

<H�v�R6I�
'6���p�[�b����	鑺N,��pZ�*㚫���{��/n{%���0��ǫ6��_2b�@۰�k��h�d�5�(���U�����4ʋ��0��9��^<�>J�W�+����
���W�,��$�?��$ �J�)�o�T\�ɹ�R�h���Yń��6�&�-����?(�h�q��2�g����I�S�6,���F�v��_9�Zq~�ڶO�/C�!��P*jK���LLA�2E��HW��/֋LX�,���$BK]0��	����\��{%`�fG75XM�}������I
#��X[�G��%S'��n0�sl�X����׀�Sܲ�I�������c5�F8�-��A��#����Q�����������������ݞ��^}ׄ�fFn�1c?ك@W�7����*=�۳�1���sf�yKvx��ߗp�I���Pay�p��W�8����eq����5Xi�ɻ���_巌MRJű�`�ҖF���!��R%�__+n"^��g�-}�SG+꨿0#�,��ˇw�t��ȕ-��g��fl)�2���X�or�A��'�-t���`Yi��Z��%���/�['A�E>�$b�ͱ��Ca�_��cΉ�
��yX���-�z�^(�ɽ!������?�m�X�,�E�z+�6���(\f�M䎔�ɑ�g�􂅲^c`=�=���~��R�~��υ�;P"����U�8c���M3Jہ��j��)!	ς�X���h!6MH``�ǩ���j�~܅��D�nn0�M��6i%��r/��ޔ^){�j!�e�ă`p.�S�6�z��33H��_g��ΐ��1r��:>���Y���MC]0(����f-����"�:遽m��K*˨|]�I+"J�/�Q�.�cO7���`�Y���O�>�6;�|vdDKl�e�R�7|<	��)P���)��ҙ�lD�Q5��������<��D�#��~�4�FV���?�b����)%|�I'	���Y��؂���ߪ��-��,�6p�c�=�y����U���b�*K��Ҋ����k�R<�3������8��O��s������ ޞR���Uad,/R��:3��r�ϟ�\���V>�P�0�6/y�.�:$jz��%�Q];P>c�1NM�:�gs�|y��E�+��K�V��NSc��T�d��q{�W	��Z�7:��`�R�+�S�c��15���dC�-��n38�`��N�	��1�Q�8��?v����-ful�.��h�)����
���-ۺ�kh�Gn̑l�k1� �_5��E�'�SY`�3�ю'�?�����O��B�$�I��nK�bϛ��.zi&��.�z2k_M�sϼ�1�nwٷShe���8ޟ'��-Vi/E$�5b�@��T�C�;	7��V����ȹE��Y Z�ѹ`u"�GD��ՕSq�Z��:gP8`f��okV�!"S�p���z4g��ӳ��|i�Н{�ozt������ ���I�H,
�Ž|��!6�V���}o��v��74��I�.��`f��XR��F#&LR$�-�֊^U����[P�?0�0[^�ѣ�A#7ҝ�vPuO`%4�>G�e9>ô0)�xUR]���-�!w��� kJF+�����ӹ�ϧ��D��<�}X��C����>���Co;����hU��
������۾)W�`h���*��rc޸��! �J��v�kZUL�>ϫ�<.��L�"G}��Q��a싯�N���/>�Z#��PYAQo�@�R��9�kf��S_�%BݺM�|OceKe���k�VQ�tt*Rɉ��b�邐�
=�e~U�*Nb7o�16���?~���(_��Y��W��<b���lLX��mD��?��DV�Z�z�u�2���H�ڭ�]L�A���Z�|��u���&�ot�^U_M�\p�j`P#�c��4ܦA��9�N�ƫ���� �?͡ܓ}�[x˴�E�t!���͠zW�+O X`%[>[�0���%Z�,�;;*ͻ}��8���������o�/?(�(Zn��#'l���ۥ�w�J�Pӣ���I��x�S83b*���LBhﴉJ�Y��\F�7�%9�~��4o�zցdE���N�SLT�<��[ �\@�e�v�	K �/r?��-h�0�	��1[�
��Iê��R�l}�i5fpv�{h|�\��T�YZB���	�یH5i�����1NB5u`SQ���U�P� ��'<�{�͹sEih=�Lr�]�Sl�a����X�R.A��Uo��'�-�{g��W+�v��)���i��_�.
�����:�'���>�Fy v8[[J����lP�������%q�.�Ü��H8��>+ԥ�������q��F'��#m�b�7��0�*��_�%_��Zob]Soe:zny[7w����j*�#8�4�4<"���L������ewHD|���Ʉ�@���Q@�-L���H�)�·�Hv��8���{2?�T�Q�c ��4#{�q�EP%+5�,��]�{�A��l���M�8�2L�y��+·b��ޫ}���<>�As�FD8 8�2]���n�)wN����sl��O�ʗ�g����Y���'`B�'��6N��h����C��
�u.:Z������1h��pԸҹ���z7��?H$�@��~�{!]���F��u��3�����~j�����
r̽��M���F/��+*Xܓ�w��9���LA�W�o��e+,�c�w�F_�mVng��]���;Ŭ�2�E1�-������\Z�m�2Br?��{>��jGU�������wx_u�}�<���GTUu�-�GJavL��:�� ^ؔ�!k��Ɐ�T���b��k�RrU������!��f����i�r<i��f���K�R�a��y���A?O���1����Ȁ�w�Mo����W��r$9+�u	L-�Ś�^>�S�b�VC�5>�~d0�\Q5�K���&�ϯ6,�0��b�ǽ�tҝ\�,f�����F��H��/[G�@�扨�}J�\;�>g�a�N�U�-1޳��w�yǉ�'�γ|[�9��?�c�Hd��!檄��d(� %G�?pV���cFH�QcI���;t�E0=� ~ۗ�pd
�����Ya�M��q1�����=\����3#�s�_�+�m��9 d/vd�ܗ/{� �$dfbEˏ�M ��fmi�k�e�c�U����0�$�ƿɭ ���<����~��_�?Rh�T�6��X��1B�u�˺N(���:~�X�c�y�]z���;��7�yk���ҸPp��ւ����6���{���p�A�j�����D�2E	�Ύ>���;j�1�wj�|v��I�� \F>2��2��|D;���l���.t��]��y��-��U�v�gYsA/�����D1���T���=t��8"G8��YZ����+�|���34�M4���\dK��L�����E�@���?R�3UY���s�1߬Dș��gNpwo@�܉e�˽�&r=1g�a��i{~L�gSj�K��!���ej�zD�h�0>� �/�6  �r-�K.�!�2�-t���%U�$�9i��x�-� h���r�F��&t��U�el�'N4����u<�Ϡ��Ó�7�����ޜ���N@m�3Mr`O��� ��;�I��\�&�' �"���^� ��uQc��b*(���X�*o:���M�E<�㞕^u��\:&0�GI[YFؘ�O�#Јz��B�g?��(����\BF}pTO�YF�q�ś���]5/aѥ��x9����^X�}�]键�Rm��3���Y����嗢IM�[Rl�	��  �mR=]M��a�d����MҬ�)��C�?���c�����7.0�kyc��:��ެu=�Q.Id>T��B����g�w�yj�o��1eK����ZyST�zT����|�X"��7��`m����SS����B�'����d�-\8�nĠ�`k0��ښD��Qˁ׺p᝛jlb-�p���A�'E���_��1�>�u�(x\C���I%k�=DK�5�������Y��E�"�n�L!��?S���b�����0Kcn|ע��#��&������2<4;���w��~|n��7S�:)�?����cȄM�i [>�&25@���z̌��a�#�v ��j�.�ư�Z �qħ"�xvK�M�Ĳ7ZZh&g��f��bo\�����k"�`�ι4ص��DEf|�L��o���t*���<� ӫInL>
7|t�B!�G���AI֧�G7�+CIEԎ��N�ȡi#t$ހ�ֻ��9����У0D��t"�#(�Y�/J�u��>4�Z�����>�7q0ڡ�U#:0���!�(��k�#+�!��d/�XB���a�-��X˅"�O���C�m���;7[�Y��y9�ײ��3W)��h� �E�r�U�䛋�\�v��U]�`>C�I��.��Zw��������]�B����M��R>?#*�P�LFoz���09Y���������������e�Qa�+擘�"<��ָ*Cۙ�K�@��[�e�"�*��P7 �26�� ?o���9;,��W짺��գ�L	�~mrY?�+�Dg����Ѓ�d9���><.L3;!��@���&���{�N������^�����hj1���ã���$�2�⋊%+�7�Uהx� k�С�;��z(xܔ?E�V�y��o.�m 	�N%,'�3g�i�Zޯ;���,����ܟW�$���0� o%(��Z6*}��l��:l(�(\��!>�uy	�-1�>�8�͇�F�WB��T�:@Y��1F{],%J�-�0�o�΁���ƈӦS�jG���[��\Q�q����Z� ǳ?~�hBh�	r��[����Z���l�1*5בFv�)!h��q��ʤ�ELYk���N�,�65��A�#qy��mF�B?Ӑf�C�Q��'���ԍ�s�����=�=�h�d�iaB�j��5��I��#�M�:5���Ԯl�8�h�v����F\�:\.�@�\z�:Z�u����W��vi�0[�F�bJΧkЉ��q��Í��HI��άO������ނ����E���a]b����Ay>*���=e���3boz�nJ��w����$X6*��,����<�c{�`�]��饊w���|
.ɵܶ�GQ�h���܄�ʣ)�z�����(`�n;?��Q����#,��I�+&�,�3<ެ$��K��'����8A���J�+��ְ�Ю}�O<�_��wHF��_8���]���C�)�xf�ȯs���4��("�ם�־����?`S�F�جK���i�C�^��&Uy�V���b� d�1��p%�Z���z�����3��~�s!]���F�`S�G�ǹUy����kI<
CK;���z��r�F`@�+l��XM��w^{��h�A_��`z�v#�唸y���&mǸЮ�.�x!�}�H2�`,�>G.�KU�ۭ[�m�H�2ӵ�?��u>�=�GF<��}��C��_�x1�&��sT�u��!G;>�L�b�����oG!ܒ�BK�T�*{������ݺ�cn��a���!v�fr�S�I�r�@�����
A���u��f)��lߨ� ���v5�q���uM�R�{6�L���d&z)-�Q���:�d�b?X�C�����e�����4�����'�$0 �b�X��atC�`���U�d�����"���y��u@��ޡJ-���:�a���N���-B���wD�0<w�DW[:.��ɜc�-d�>�����(�|Gc�tp�����c��bgصz�t���=B�x~l<�pAӕ��3��qa��'ʢX����=�|�xs������y��~!$�j��/�2E���{��]$��E��>i���i��i��E��"9���e$�`L�~�ж�����G~�	ߐ����k}6�A#�ɘQBh��˫y!�Y~�cm�^�u���{��~�y<����^bP����?�P����4v�~&E�tm�y�j�����~2v�."��jrݹw��v�ɧ:.w mRe2&;��X�D>�'�l��Dm���r��@�ںZц<xǡ�Y� �Rz���;�1�#EK�N�!�i�'G��.Yˤ-�9��+�(��T�3%�4�H����M��b��(��@f���*�3F�I��~�b�D��}[bN(�@D��e��r���1x���љ{�e�ؖ��������ޔ�O�k�h�B�Q5���Ϭ�Q�K�b1���3EZ�� �� ��9���xG�U�q傌���5l̙�OR�Fube}�&Nehۯ��P�@��\�_�8~���v��Ĕ�Nq��3�� `���2������IUW��� 93�-�`�Q{�u�������v�����:�I��^X^m����4�uJK:��G�F�x�O�+Й���\(g�W,�o}��C�\�ٟ}Au�O��=Tׂ���7\)o	��6��\-���4���u��������~)&��n�tU�9�z}0�hfCK������^��ȍx��^��ZN�	"Y���|�VUi�����w�V�F3�P5�V[��O��#�j���K�/�ݢ�آ�㯑�"�-���a�8��j��;�p�|~�:�[�r�D�c췃P����&	��H��Α�s�RQLĔM�i0]�V�)�5*1��|{o�{Ȍ��4cg����k1xUlA�����hC0ˠvO���x���.��k
�(�ZW<�i�|`�E����(��xR�����a
�W[i{<�#����`E��
��-�"�
�7���/�sXU7����sh׃VK:,b�YM�ŝ��$��qtA�hD����[��K�,l>x��hx��K��?7��Z�����@g�>c���&_8Jf��jK�ԧE��Ak/�s�x´�����c����s��+c�X�%�%0����2���j�g���!Br� Kѱ� :'%�&��-|�7g���`�t��z2�5�C��8�Q�Y�;���[�-��R	z#_���;���ͤ�n�d���X��-&�i㳜�2��e����4%�n�B;S������៲A��A�,i]�Ȼ#�@�Ǚ���i�*���^֓zC�'D��#&�Z�J�"!�(�:�A
�Zw��g�ĵf�0�oYu@�i}W"��r��6�4U:l�aYi|׫j����o�ot�ˊ�k� ��mI���
7 |1�.!d��D��+iN���7b�0I��q���<��%K�#֦${�������o�I!5�O0�"	���5#%j���u���4��T�S�>�0���U����Ӭ!%%���7kxM>��s3D�����52>�*��Xh�6���>� ���>�;T�=�����ׯh�ܭ��)�w�h�DN��r��X��xF�v�;MU��j>�R��j���c���;��K�"":􋝤Q�1��>|��#_PGfMo�p���F9��"��?�k���(�x���e9�4�H�Ϙv���L�R*@v�����W�c�8�el�P*��[7��6�P?l�=��d���v�Wɬ|Plأ��[L�G�mr�?���D{L����`X��0�[�ML�[0��64��<��8�������.]�7^(,��Nwj���󖴌�W�+�o�ˋg�8��$ױ�� (���
�y�w��xy�Ehl�<o͎-K�� ��%���	~���Z��;i� ͩF��� ��ߞ_F�g�(���Zs޿� �luc���e����~��rϬ�I��{��8a����1B�i����Y�*�Fx�Q%�r���o�ɁRƥ��S����j2�[ ��\�ӗ7�7�" ��F?<c�h���	�m�[ɞ���Ԋ�O��l���5T�v��Hh�ʏ�5x��B�vY"��N���	55W��@�K����	?E�JJ�'j���
�Os��uyW=�O|[�aZ�Ѳ�@3�@��ow��U�i3=�uYv�;^�#.�r.�&��$�:�{�������v�&[xX�ߍE�6m�F�q��ÊhH�������-���ޟ~д���Q]�b�-��޿�*��4}ٝt�4b�o�j�n��Ew������*۞�b�r<.��}ć�tzV��%.w�Y|���������6Q.`���V��)*���h���VE�MO�?았Q��֖:y�#��}�sx�+#�,k�O���p�(���xC�`(8��
٧Wf+��\�D��}6�f<l��/�;F��8T�Q]����@)%�͒XUs���J�E=��ZM�ld���`�,ӒBd���䤅AGC�F���@$D����yw�_1֐p�o���5z�����x�n[�~��]���F��$0�ҫ��,�"�(9
��Г���Q��F��+I�wX�\/w{ʐ�%@�A����]P������tfmDE���JϠc��ځ_2����)H���#ۊY�m�t2��?R�F> �GCH�Ȏ����ֵ_�ik�O�2@�T�l�ub�G8�LD� �)���!Y�}�_�:Tu��"����g�� 8׮T^�ͅ(!��df����ל6r<���W��WW���m�٘�gڷ���(���@O��n�o�Q�]M�)��9:�ɝW�S��-G���P��6ib|fC�2�l���
�j��υ�T���$,?0�-b\8���9t��35Q&����L����%�:����@�zF����JJOt���)aGXN�q-�wb ��w�6�����a=�[�m�H�c�r�dn#�T���o�(u�KG��3p�J|5 c�}����!�X�t՞�=��V~��2p����#�T�a�Qc�ߪ���c!=JRy����1�8}va���NʧX/�YQ܅�B{�$�t�E�k�;b���i d���Y�CRo���a$Tc���*Q���<�-H~#!�m�M�B�56�-�Æ�B��i˨�}̤�?~W
ccJ����!��4��;��y�T���^�P�pD�I�-���$��曬�1�0�o�?j�nɞ)2��"�	����rj�0�w�h�vMXR7�s 
��2c䵗��jD����9V���n�G[�w�������kYa>�og��k�~1�PB�-��Z榙�Gf+�YH�VU�+�&���y3"h�4Kɾ��i��* )��+E|j@#+��m�3C񆸬v]��r�D����@N|L@we,���`�17m��?�{��:U������ߏ��_�h@)hh�Y��n��d� �`p�K�P����>�C��.m�k9�	?x$���c/��>$��יTF��C7�e�,N����ή�����yT���	H���x�a�N�ƅ3{�6`=O�Oܨz�3I�g���� �Ժ�j�۬.r�u?���@ܷ�X��:���@�����̸�u�I<:�ֽG��>F��O
*Z�6ȧ*F�gmhMv�����I\�`}��kO��Tt��Z�����)�b	�S>\�>-9y���B͸q����)�9nˤ��Rzځe�j�϶��;>�
,��ɁJB�p�ff�V�m�RU��K�9���/s�0��x5�����&�R��j�J,K]������֯NOm�����8u�j5���K|�ы��{�/���
鯷��ؼ��	N�Hu�_�Y�2Rn���Q��i��_V�$5����J�笑�\u�Yc$�
���k.>l����
lnb0HbvO��xy����zk����ѽQ��|��qEw��E�]x@�V;
�<li�i�`,t�]E-8p
ٚoV){���#��Ұ]r7�p���J�s�,8�M���,/$1'q�3x�E~��6mZ��p�,)��QI#��R�E��4:g��V��	^>�����J�z�g��Dε���k*����`���� mӁnI�(��XF+�%m���wܨ�����$���,�~cr���N;�:d˞Δ�����r�����~�Z��O�B��:�ݓ�&�LV���ؼ�~.�3\���Y/�7�ل�6�a�a���"�%Δp[�9�&�&��4����QOЎ�a��ͦb;�3Ώ��d�;'�<f'� [\ّ]H8���#��;�o��I���HLpa����V:�H�g~mj�C��9�B���r������ڝ|��6c��?��>p�yb��*���z�+�S%��M����Q������A��60�A]�]b��'%j�*'���2Rm�bV۰�h��ɘ�������;lW/�*k�a-V�P�;���h�]؇�Y���lQ����(3q��nW��!�}*���\E��h�����B�Ŧ�Z�
��v��UW}��mB��O��N�W�����n
��to'�	q���(vd�n��GWƷf\�6�{��V��1o���7��dO	?�|�{y��`}e��O�q�]1��=vw����h}��P��L�2���� Н9�A�����|�-�$��|�]_=������&�8U��'=���V!	� 7rY�S��$��F�"|L��&����\���@=O�r��A���o�&K/#]���<65�Z��(�����G�P���3�Z����bq��^��6=��~&±'��F&�3�ީ^fkAZ���vys�w~t>�U&&�:�
�8��W�D���!�&;sx����2�:�S���DMe����Cq�<9ťϽd ��q�6���-��DM Z+���3մ)'�u6��ک#�?��&�K�ˋ/׼4\�-Uū�'��s,�i�y2ƒ��`a�c�<��4�ٷ=���MQ�=�L��%�)W9FL�\�0�R���������S��Q�s��]���߿b�U���݉�=��_g`^��-����!�*$�c%��I�|�zY�5��;gB�$#�=ɵ�fzg����욆iWn��jj"B��ԧpjT��s�q�c����A0����Δ����5 X�i���*g9�eb�A�. ��lJ�(� W*� i�\h�^Kl;�ݻ��c�C�	0Dۤ9�\������6&�']�	P=���"C!H��L�ʕA��T��`�O^F SP+��u�/�|�A�����+��a��m�1�ɏ��m]��f1Wx(�E�P�(i�3���u[$��m8%.�N�K���I���8�ф��`�M׼��P�au�"�^������cK6���_��"��Q�9�Z�Q��^�ZC��p�g��zҸ���Yn���R�0�a��l�?�r?��T+Ƙ1���ۏ�$��J���9�\B� Q��X�Jl�WQ�V�f�_hi��V�aL��w��>$\|��F�elZ����S�_�;Gd�'��2���XL9⏭��gl���5��2����z+�O q'+g�9���~ӕ"�v;�� �!�8�F�S�I�Ϣ}� #���[r �����]��yy�e�B${��:9.[�h ڜ�E!����_��(�z?gq[���U������Hv��u�ٲ�H�j�z�@eߩ��Ap�+�LF�9��V2��N���*��f�XI���&6b�Y�k�y��ft/�Eg�.�e:��s��^e��5n�sN[b�#{�l|�P.w٨`e�@�7_�l����)�{�J �������dEU�)Ȗ��ՈY����K���y�+C�2�~�qaU�׮1-�'���&�/�����7�y[G����M��ԩ<���]��/��4!�+���o�y��	���pQ�<��/�('�%PҭE)��6x����d	��+N>��m%,Z��&㵿��T�
�{`�v�˅Ǧ����xㆹ�hfG�5�Z��ۀ �����/r��H/�ju��I��~>�J�4�+B$ ��#P���L�������]������J�կ�xq\\�f�M��H���?�l�Qi-������'�(�Qq� g2�pO�JiI���6G�x���Q�0_t?Tq��J��C�tO��K�0L���������I�K/�*7X2���_nPKx��Є=��z�\4x�%��cfB��X�@ }�� ��/�I� �i7����%�(�굣7��@��/���7��p���Ӹӣ�đDc0�Dx7�-\����e�^�@Qz��*Xkٷ����WEb���J�����}RU�f�%��l>X����C����B*���8㫴1�0f�qK��x6N��k���=aa4=���Z�8h֛0��깍�p�����wW,�r��R+8j��'�w��2�֍���R �D_�D�^���g�P��CY�4�k*L,7��˂9t������gd"l�Cg������GAE@Х�t�����Z�倊{�� �/�x+A�
Ɔ�l$=�T�W"wH���d8س������u�H(q=�x���UϠh�m���,5y���r6���(�|M�������P�`�(cS�C�����77ǭ]�����ϠyP�X��`��s�-�La�3E_K�&n���Cϝ��Z��!��`���Bֺjz������znK�M�h6D	_���H�yۅ9{K�4� "C�{�}��x76�	R�Ha|�g���8�1-%���A	��)�ܒ+���]�Db�;��fF�;"-�8���0q�㝟]vѾ"E]�/E,�.Q�^7����l��k"O��j��-��w�ED�q�eQJ7��<��j������r��Ҕ��DH���S(��,Y��-S���%���ϕYV����i�b]qc�Dç�Ĉ��{�򄀰�IW��Q��o�V�Q~5띿p^!=�B	��g����j������Hꘊ�Y|��b}R��3�hŃ�݊�镗LP�E.��3� � aR稰��"�dǣH�Ҭ�:�-��� ������g�O0��y�o:=Y�X�Q�/>~��&k">g��
y�ُ�&i�KZ���	S~�;T+���X��PL675�m`��ES�n$ج����?�d~�-�>n.lj`i���H�',Q5�&�_ۛT�O-o�)~G��i���v %r������i-W��,c�k,���h5z�����rY;-�������ig��L��?�+��n&s���4e��F7&	}��D�2&�,�'���nRn1S��W�ip��Q��.��i���P�B@k6�/*��vD�������������[Z*7����5"�2�5���~`ZĹhg�Ff~o�x5�6��".$���R4YӮ`�|Ĝҝ6�.o#P,t����~
K �."I�,>
�|$�!�q�����-�Qq�7o�sIo}�[��)�}��Ӫ#Ap�$H�Q�e���#����	U:l0����^��#R�*��hu*�24߻�� ^j>{�0�R�U ��("!��܊qSk�λ�Ka��<|�����q�W�CX58Ɗ����-�ǜG>�;���v�c����v��z�)2�Oh�?���a\r^���EZ;� �v'EU��_>�1�w�q����+P�8��0��l��bz>�9�#�1P�|2o������9C�V���Z8گݕGq��e�覕��cZ��X�*m��x���q��ESeg�*I��7ʶ6wd�?�������4U[W�X���O���L���m��??�[D�<ԑU�!�m|�c0�ڨ�KL�E��^+�#V]��}����Y
Ǧ^Px��>ja��êQ�$`���ۦ�t�z�ai���i� ���/��xF+=Eq�� �5�;���g� ��|%e�6.��n�}Z�;v+��V
�3�D�杞�zЧJ��(��|Z�C��:�l"�}�w��Ҙ������������R8n���p8oBc�^��^Y~�'F���%��t�Doا�����@S����K[-ʁ\�l�@{\�D@� ?o2?�+�h�	\}�[��M��������l��h5�Wv
�Xhr9���ė�o�VY�Ŝ»��ۈ5�������*[0T6l א�j���;�'w�ԷM�s�@b"2=��~���΅�a�e	���������,\����ž���]�ҏ�v_�p�0��d��.�L��:D��k���(	v�Y[����.r���-�3��q�N�÷��H��xx�\��kc�6���1�С����8b:��Q�*_�>'��!��bX��o�$.n4�hw��P���t*��?�o�0<����q��a�ߥtZ�w" Y|t�u�_���v�Q�tA(mx�C��)����`_�޺q�?��Q:<�� �#�W�� 'J+P-e,84�V2��5�C�IG���8����4C\+� ��}�#f<yl��!�F?�8AyS]k���2��)�u�r��s�\��h�ʒ�k�Gt�֨����,�`�)0���`��Et�2'�C����E0�\A�n�䊌�1CD6p�t�8��z2m�욊}��:'~���]_��F���1�Kx�yz�N�
-�b�	���/TF
�+V(�XwYZw�\�]AI����S���>���hZm�}��9�P���g�2�Kԑ������ۗn�m��T2=+�??�/>���Gp�	�[�C���_�������T�u�rfGe=`LG`��O/���!H�TSTba�����
g���4��܍��Q!5��f�g��ĉsrɖZ�2���t���-_��%���|�$���I��g���|MJ������v%�41/��@-�S���y�Α,b��C��;��ؚW"᧦�˦�ܳ�Q�0j��b�**���gtm&*�����S��;ܯ..��QmZ��@ x�C��J��'���KaԽ�N���-�J!m� w��A�Z��ή�[�p����c�|Md;s�Q�����("��G��p����5�ce���e���EQt���=lU�~�_�p��j��f�c0ae���L.���6\#O���#�j��כJ[��+�����f2�`�w���0������7���DJ�� ��\a,J����Q��$�?��[g��3K��w(��q���2p�Τ��I��
6�I+�W
�u+_�t�q���ǥCB�$��H8KD�L����_o�5�SNĐ/v"Xw���D�K���Щm�?��\���% �=f�mX�}�<j�f�wI���.�U��u%���ZE��������R���z��^D8-�Ė�9c�!����-A7���T���Q?Z���v�ټn��:�:������]�+}w�f������"�#���d9�A,*��%��}��V��fFT�K:px;�=��g�^�9a0�^��88S���.�aȀ���o�i�w��v��W��R�<�� ��r����<C��F�R�y�_��L^��]g�����-��c^�1#,<�O�'��t\����!�g��lɂ�R��!NAJi�u��t.U� X�_~���Ν�/:�&A�h'����n�9��OYm���)F+�fh�������H(�l;�]`�0��6�mf��,�� ��6\�K(���M�m��iD���%��c������7���+��lƱ�x�%�^P�@G�%�Z��1��Q�3����k5���?!�"�t�!�g+` 7�G=�jC�%���?�n�b�MD�[6	ࣗ>(�~w[�V��{�u����� ���_�6}��'��HfM�g���}�t1�q�~աS�B�g]�J1��c���� #�"��'�]4��H���H�]{�"���/�<!.6��77i� S��0*)OQ�F�֝�-0D��e61�7�$<����*_�`X�����9>UD�|(�8k0ֱ��R����s��ZMb�o�VYǽ���<bB�M�����m��@���WGX}�A����<�6���"� p�J=M�!�Z����Н�L`��U�-l8�,�#�R�\y3IU�ňu����ꗑ�*Ś���� �R���9��d�Q��_��}g��_���}�<0�,��01%�y��':Ā.�d*Q�yd>�Ѵk0u�gx�y���ˁ K������HSN<TPk�tL���7�Q]�7���`\}�˅�SD�=����h|Nd�ݓ-���n�.�`Z������5$CQZ�ߐ���	-�
��Z��b���7�#����뺗&��VS�1O�k�	�:j�5_Q_Q�C�`Y IB�q=��������yJ�1��ĸ����Fn���;^*�Μ�&��ͳ�/F2����嗼&��ntgSTN�n�ޟ�=4�s�iσݻ�t�@�l��$��ۗ����WօHW�Y�k�8�Z�qk� |O"S"�����s&ZiO�g�b]fc�ohH�[�]"�B�Z�{46��S�n|	\�:�o��dt����C�> "A�I���
)\�|cX�!����""�V��@=7ԟ�It͎ �gnc!����#�~$m���*�軈;�������0���C�6#פ2���u�Z94D���\>�9V0��HU��]��!�͊6�Tk�4��PI��s�&�G�Χ�����XZ,��X����L��;FD��H�H���aYpܟ�s)�\�hB������r5��L��:Dv���U�e?>�I���S������=Q�}?����O�~�#@^>��Q#y��P��yo������9(*�H�']�Z���^�e�G��:�E��`%����*�Pʉ�C��ݨӪ��eؕ*�8I7}66\�{?���ȅ����EW;��@U��sL�ϫm�+.?�D�m��S/�Ҋ�hW�M�@L"���n^ި+�*uB��@gU�W�y^�����j /K�H5��I;v��i��세f��ףOt Zjԡ|j�)��xk[�E6��e��@�="� ��%�\���"��N8ZMG;ۍ)�[����(W�Fj���ŧϝL(���Z��*�S2{l'��{���#��1��$珬�(���f�8�s�uQ�B��)�Yc��F*
�%�#x9�Ro=ɳ�hXƗ�]S����P�[���\�Eay���\ D��?.vh1	A��[{A��)]����lP5|(v�Y@h�w��:P���Y�HJ�i�{��5	�F�2@�lA����V��B<���'܍�Լo#s�;���=mkh.P���a�7 �C}��p�2�i�����z(�����3v$wkו���iBe.���K��:)�4Ëq����v�s}[�K$���s�(�g�x�4qu-��<S"H�e=9��E5�;Hޑ�P��q����b�������*$S#���&�b� o%�n��w����ж*L^��Ԅ@<�E�o�u��F�Yx�w���|��)�$f%$�GQ�	͢焈s)�A�}�|��߅��?^#Q?/�,+#�Ӣ�n�+�q�,]	;���Ú���NF-��K80����z+n��6�5}h��<޳��U)F�n\8��]Pp�ʷ�Z)�$�75�s9�ѭ�7e`׌23֍X߃��`���G1v�<�4�7őC�@@�y���ߐ��䯵�1��pt�.�=��zנ��2y���~N�[]�,CFK�~���c��S�!��Zk1
�ԓ�3@�COF��Z+�X�X|��wm:�W�bA.������9��-�m�[���Š����L�2A8u�����Ԫ���m�_�2�6?�5�>r��G�.}Ȁj+��1�_�B�a�$&	T�u���G꓋L6n��[[��4�K!(��Q�BT�Ǿ����rY�����݆?�j!:��f�ne�	e�r��{��V�������T��KP`��0߷W��tW��oN� �G�C�;M�}_C��{�+����-�s��:v���b��EC]d�g@���E������_P��~20���b���]N�tr@'#3�D�mݾ�+���Ѵ,vb@ezy�H�~J<�d���.a�jNA��-��2��wW���_
��S�E[)D�ں��cQ{jd`B��6�K�('��Gr�p����c�{��ֵ��mtG��=qC�~{�pU���R��˻a�����-�e=��F��Û���( �����:w/�V�7|�{���$��Ekn�Q�m�iRFT��R�������C$����Mֶb�l�Pt~Mz��� l���6���ø��B7�m�ZA�̖��~�s�c�A2���@��h��m��yM�˓ePuv=Yܟ������捲L�c{��D�j}eɐ�{2�c�n=@�Ibsj��w
?�v����q �l�2���>SDm�"�{��3yg���^�j�i������{2YXa�`��ƨ1R���������\�G�T�Y�f1�H�V+�2�#^�3�H4=� ��>D˜{���7��@UI���Ѝ3�cs��?؅�Y�Dhh����Nn@3��e�����dP1�Қ(9{�r���볠��W}�c$���8hZ\��y
��R�ZK�����$��W9쯪\9	'�x��2���d�����$���r���eN��5�@���o�k���'����꛽1�SƢN�'3�` `��A���%I$8�Ƴu ��$��{��+nu��	��J�rx����:�����"��Q�>ėu4û:Ɔ,G酃FxjO�,��(!�\�@g��P(�/����\���}s�O9L�Tf0`��c,���.)� ��Eq"\����f�ͪn�?j&�)Ui�n����7szL�O�#�{��3n���� ȼ���ylt�ѱ�"���{U�z�I�Eݦ�e��"��5g�g��(DM�j�>K��	�щt�!���i���m��SO8g*Bjg��W	|�I��S��a��|���2�7��% 	���H����R`�ă�3i��VH�	5�����a�⑪�h��j�cV�S��Gk�'lЀ��ޭ�0��[O�cCx����0Nk��?��1���|a��E�6φ7m�xA���sP�
C��i
8Ғi����E߉�
�"X��"���O�[�����G7@�5䢔��e�8,Q�.MY7��c$#*�q�z��C���y�Ꜿ,[����9l�����7�b�f������o�>r���Q�J5H�u��6u3�*��k~Ux��+I� u��R;I��y����X8�V%�Q���Y��a���y����w�QrL�7�@��:�t�@d �\c8r�+=�Ш~U�8�@�'4�":Θ���QL)9�wԔ�.�����u2A�)�_ٶ�!���a6��"�=���q�9��&[�}&h��!�OBTa�Sx�T%{3E���Q��;�#<�o�͑�ӎ(� �`P�M�Hj-��7@;l�r��+��*�jL��:gMjV,W�Hгrm܊����9�yP�	�5� ��J�`ڏ�o��1�)����p�)R3a���ݦS�V��\fbI:�����A�;瀨�D�󪬊OfJ�Y�¡����	�m��VM&��Lp�J_���I��D�qJ���n�S�QV᭲;� hR�߇�O��tQ
p�m�(%S��%�m�Jw�}܆d�N���? ��8��B�Rt��|t
�B��p�*}�"�B��rO>��Nn*{Ws����ɒ
�xo���#����F�d�JN���WxhK\�԰�������81!�)�)�hd��	���-���R����@+1`Ծvi������ڃ�f%�
/��d���Х�O&��^���K�@�ùc]��#�9��	P&�Y�=�Ϫ�	�/r@F�S1k��tH�����]e�"҆��<7@/0'r0�8�A�F����#O���n~�*����Eu��V�X�PYG��X�Zt����_q5�V^?@�=��&��ʇ[�-��Rޛvks���Fi,s_��t0!�&X��`�n8��W��P��!Ck*s�J�����l k�kEMv���2�nɰ�AT���qz1�����a�^M��b��=��G�''fl�V'�ێ=?Z����ئ�!��4���U7��';$K,��ydCo�Y���5T�.L�4 Ix�)�y��5y�?��o0��C�2�z�F>3��b��R#����,B��"����s0�����Q�T���'���n���`Pų-����#!���k��UD��-F?�h z����"�B7��#�ֵ_@�zY�����r��+H���#\ۥB������T�<~�c���6��VՏD���ى�g�� �,ciI�*Y҄���JA���.�<^�	�Z�W�A�i@�g�P�];�!޺o.C�"�D�Ӏ�����p���GT'OSPoi��;�!C���>��sTL�V�^8J�P]�u
q�ⴸHA��ժ�@`��p}R��#���	����� �x`u���Lۇ༘��[�"�N%��6��e5�z�I���c�6�����u�b�����u�k�^���dc��G�ӆf����",N$��9��C�^�ӹC!��p�5H���ĸ&�2Y�����0�ND��H���0���s�ƊGƸ���ݖ	J����S��?�G�
�eJ^�W�nVTs_���H�(~�dwCq�$�a�8�l��؍�Q�_�Gd�z ������?*9�eH��t]l֋7�c!�����	Ɓ�'���9[+~��ђ��X�b��*Ļƅ�_�A.P����� N$���
J�඘kR�e:ƻ$�a�����   �   Ĵ���	��Z�T�
0Q�ȸ�D�LDr�D��e�2Tx��ƕ	#��4U�h���ƦE�4W�Y�4$�P�\���L��/˼P`��i��6M��Iz���'���x�e��<����6��p�T�5����G5�ɹP�8'�i
�x�weQ�u���%%�E�jh	�O qzcJ���MAT��!PN_�Sj$_�|�q��45�����ҡ���ѧE]�f_�-@�V����U lۅ�kݑ��O04���Ԯ0�� ��E�&^��`�#�P��27�ʶ��$	, �|Q�q�iY��+v�m��_?���ۥ<��t0 h�!��	Ҡ��q?���M`�U%�d��BR�LUQ6����@Ӵ��}��o՞(�R92g��b2I��i��r�B(Y���F�EyH�X�Nڭ{P̍��K)[WV5���\�)�ܒT�T�`��s攰�2���j�f˖��(�'%�T��O7J��S�����}�A�'�֌�撟���'�\(�� +�'"X��`��p��qD��O`j���,������<	v�H����<A�.�~R�#f��0��ϫ]@��!����MT<O�� 2B'?�8O���@-?i\cŸ\x5,�,qs�m��d��`�L9U�0�G�IF�O2 +E

=Z���é$,��jq�0�Op����D��?���-w�44��%�i���/L�#<y�b?�3aT��L�� Y�%��)4��G��O�M<�R�ȟ(�p�
�k΍0��2u�T(;�)-uT5�p�5>�|� ��ǘZ���� hU���Q�SL�)���:$�K쟐XC��s�dA"�	��/	V4hw��<��ęY�D$�hk"mE�Y��OV(��.R�Y�r�@�ш!�i��g�.*n)�7�|R���Gxh��y�g�/syܵ)pS>:nR�)Y�C��d��"O� �  �                                                                                                                                                                                                                                                                                                                                   �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  ��   D  �  �  �  +  �6  �A  @J  �U  �a  #h  tn  �t  {  H�  ��  ύ  �  g�  ��  �  ,�  n�  ��  ��  9�  ��  ��  E�  ��  ��  ��  
�  � �
 � � . �"  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��	Ty^�� Ui3n�>>��L���$v�������`0l�S�`R7P��%%�s�a|b�|B�Y5$���Ӧ�?Cg��iЈ���y���(uY����6�l�c� ���'1d�F{J?9�e�¨a��Y�>X�y@��-D��挚�n6~%���)#/΍
s�*���<a��@+A�n��C�)X^��ĉH�<QЩ��$+04A#B6v���$fz�<A$+�% ��U²J�3�|H�� K�'6�I^�O��\IE)��,� �cʁ�z�	�'�f���W6`D@�JG�����=y��<�}"�R�@)!��j.�Ŋ�F5=b$�	ũ$D��	SL��rOz�Kf&�|.�H��`�$�I��HO>9�@�F6PWN݂��>����!?�O�O�m�Ǥ�?ZdX���^(�����5|O� j��Ql����U�j�pIB�	f����C-(h©���ɒvɦ-��<,�d0�OX�J�
|�A0��'o$|��'A�<��%e��a�%D���J�0�L3�C�	�)��	�gџ.o@p��+ȣT��O�듇�'oqOve��L;�����&&np��"O(f�ݩw�ؽXeC@�����Dd�F��Dq���w�[5	�`����!`a~��n��kܨd��aKϘHv��[���
2]!�Ͷy�X �kZ�7��X�(H<
{���G{����k �ɢ�p�VH	�}v�4�U"O���BF\���%hX�bD�x5S���'剧�3?��ݒJT@��E��lZ�T1AAQ�<y���3��|��Yc�څ�n�W�d?�O<hhƋL3z�8�	�_=,���"O� 4D�A�<!bPc�@�+
��f"O� z�NX�|�<�D,�U�X�$%LO�8珓a��<RLW)b�"OZxj��B3'R�Q����38&����"O8`�	�e���۠�A�w�m�"O�M�g*r�"M2F��l !�"OP1,	��T��"^�Bk����"O�0@��)5���{�@�C�8��"O��Q�i�6��U�O�TV�Æ"Ox�ǭ�m(<2wn�g@�hq"O�8VfN 8�f �[�"L��"O�<b�(�[��c�K�bt��"ORĳf�N>qC++P(�����K�K�<�O�IԬ���`O%�^ЫA�K�<��MPT"�c�F���{4��H�<�!Ľk���S�C��hA��P���o�<�FG�s	�Mْ�-Q)�l���]j�<Q��5yd��b�)P_�0�A�i�<�"� A�r����
r�b���Ŋg8�����a$ڼb���(�.�(W�P2#C=D����T,8����%W��q�'<D����&5��%h7c����	c�C5D��K4NȎm*��9��)(j̱B�5D�(SJ�I�A�B�T� �e>D��É�>����҂ʅ��a�`f�\G{���U8CG�cR��.�@9{R�?P!��fV ��Ĩ���0@�r��>E�!�d�
�ECwM)���&$W>v!�Q�����U(��#��|�!�$�?_�p����~��Y�㛃{�!�D���bA��O�1IǘzU�	�!�$�8z��0e��d}�P$�	�bO|���JtL�pjD,E�Z<��'&(OHq��a�p�����0� �"O"�WG�g�ơJ�\36�\C��t����K=�wa�24Q4���n�!���p��3-�
K �Ä�o�!��K.V�Lx�-7��s�kJ>av!�D�6� ��aG�GXAǭ!!f!��2`���%�ZqcCmN�Q�a{R�$�<*��h��B��5���.�!��w��7�r�`���+�2V��Q�'E�F됻6D��0�?e��+R���?q���S2[l$���ڨ}����s�L�U�L���`���Kũ��V�qL�K�h��?���$7`ӊCP�S�q�8�j�'�Ha}��>��B���0��7D��LClx� Ex�&o����?h5^��`�(OL�=�O5��5��=i���9�E�:.D�����	<v@�C��V	$�Z�Ç�3��C�z4m��/�6�PH[�#G�(���<��O��=��,�!k5���b&��s�8��{}R�'��8SEܕ>A�p��H�M]J}����&'\���0"��9��>o��E2��>I��T�^D�����N�5�pPc2��,�y�f]�E�l�`�^�D�����C���'3`�à���tkC�>]���>*[ ia⁸�y�I�D<��S�h\&��v	�0�hO���dY	)����QGB@T�����/l��f
O �p�ƹb�`c��R�t����O ��d1�� �5N̛IL`y�]h�a}�ƉBy�Fܷ=����W"H�B�Jܜ�yruǞa�QK%@,��!ݐ�O."�����∀��@�9Ҧ��ac�r�<� �� L�"R&����K�[�&� 曟PD{��	�u�܄� �f�tq�M*@O8��n�
u4���l˺^�q��i �<�Oұ���.Ӄ[q����B�V��:��R��yb��W Ͱ��_$S0����E,[��$���'��Sn��f�A3#M��R���l�9iY����{y�U�0f���<;&�#x��;��2D��vo��2�{��ߙ~o��Ra�/�d{���f�Oq����\,6	0aק
ԙۆ""�y�"��_�z���҃1P�9[����~��)�'_��0��CZP������s��9�ē̔��C�(d�쭸��G.Q��M�SH<�F)G�.8h��L�_�	tɐq��$�?�6��<l����D�S�T�hݨ!��p�<1�
�1Y�Ԙ�:)|���k?Y�{��O��ػRĂ$�E@-ęT��x�ʓm�r�s��ʴS���y�ئ4���O��OV�=�өt���sFY�S*�8�e䔈5���d� ��O�QYW*Gh�0q�(���?	���g����'ˏ5�H�N�-C!�D�� ��$ƕ
L6��#䝼xT1O<���%|��l��)�/l�*S���!򄚚3����p��"��cS-V'^a!�A��6�
�4 m���_�!�$T��J�j@&�7�"8lC�{q!�dV+Rx�SD[�b��������nY�t�7�0]�f��
�7޴!*D��aG��+�0��E�[�V��L@d�'D����@�F��� fٚo���IW&\O�c���3�9��d�(B��PhE$�<�!�dǯHÌ<Q�	5J�n	[���T!�D��kS��1T��l�A�cB�	H!���,=��#P!(<�<*�bO�K !���c�|yC*n,.i(qk�My!�����xP1��9.��[��v@!�$� �<�c�I�M�|E@f��?>�!��ۊV!~%�Q�%)��-��D�!�ܣ.q6����'� �q�ɀ�b�!�� `���-�H���aC�DT!�I��qAv6�إ�q��i!�$�P2$��s��j�L00�@�
+!�䗠/.e�p(@8O��w��~!�d7T\��R 䌹���c"!�$x/ Q�b�R� �0����!�D¿:p�Q��OQ�lx(��&V�!��F�%$�e��$�Dk�b&��*!��=XF����V0NXx��Gl�!򤑝*ļ�����[�`i��UZ!�"&� S@��z�p@�$]�9�!�䅭D8�����$bʼi��L;\�!�$O04��py3�_�Gbn�0��P�!��3Y
����3RQ����f�!��#���T�,"/X���.g�!򤅃>(�г LX/$!$�(�*ћ9T!�B�1�J�
2�\	gOɂX5!��9 5���E	��Q�T�Fm
t!�DO�0��u12L/#t@!�6��#!�N&U`иr��6��8Kƈ��!򄚀sx�)����5}J�[�g���!��%LL����P�d����؍j�!���9�epu-�VHS3��-,�!򄗔X��d���H\����!�' �!򤝓WJ����l��1���˧b�9x!�$E���xh��J,=��9�ʒ):�!�� 8���㙠;�8a���3���(1"O��yt�H�C�l�sR�,G��9�"O�y��GH72�0)�օզ9�֘��L�LA1#T�.�Q��·e�d���o�2cfۣz$��G�%���	��I���Ɵ��	�����ßx�I8G�5�S�-/��uK0b�2!��ן|�I�,�I؟������Iޟ��Ie� Ӈ���k�ā0E�	�T��Iៜ��̟<��՟��	�l��֟��	:$Zڶ$E�-�t`�O
�~&��I����IΟ��Iߟ���͟��	ҟ���)O���[��I�&:J�0�����p�	����	Ɵ��	������������ɬQan��fk�#�
��O�ঙ�IП�Iҟ �	�������ɟx��Kv�0��A�,�XU�x8B��� ��۟��I����I۟�Iɟ8��)
e֌ԥ��H�X�3�W	g!����ß�I۟��������џ,��ş��Ɇ^[ڴs1K��<� ��7�Y$p��Iҟ����P�I˟0��۟��柀��Zb��vjI D�2�!�E�]�2Y���p�Iڟ �Iԟ���ş����p�I.%�����4$��Q��ŒJ���IП���ҟ8����IΟ�IП(��S]21���Es��hRI'HL��ԟ��I̟d�	՟X��Ο����d�InoZ���C�:�s"�5X^NE������I�L��ş�����y�4�?��c8��G+��j?��)�Q��8!V����gy���O��l�+:���C�G�� y��Ќ*�����/1?�!�i2�O�9O|���7���� J�7P ���g�Z-8�$�O�m�!~�L���$����OE�x!c	����:hs��H̓�?+O"�}RG-��r��(��%_�8�"!��m�V�L���'��F�lz��cq�O4@�xP����+��I�%���D���<��O1�ڭ2v�\�IZwb�P�A��D�8I熉�4����<A��'o�<E{�O ���R�(0"���d���Ç�yQ��'��8޴9��`�<�ǃ�X �y���8b��8B��_���'����?y���ybU�а5H� H74I��$Y$8���ÄG#?��6��Ʉ)�P�'6��ϐ�?�%��FVEJG�DCl(�h����<a�S��yRM^�����'���4
�nQ��yB�|�^p;����z޴�����g�Rw��PG1F���O1�yr�'u2�'P$��i����|�C�O�J��x����5��51�LA��zy�O3��'�B�'��g<$bvm�.m��MK(3{剹�M����?���?�N~���\+��y�G@����1�P�R��QfQ���	֟�&�b>UY�#KF��F�(a�f�����d�1�A/?���b�d�������/lT8�����(���nY	
sa|Rs�� "G�O����+�"I��ڸlr��E'�O��m�d�P�Iퟤ��ޟĨ"���\���Ŗ�d�x�q�b�?��am�d~Rǝ�1%�����䧚�;7��d!�fbQ'EB��K_�<i	�z�:,�N�1�1�6��1������?!�rs�fŝ���Iæ�'�@8���^��-��D\�RA ��D�I�d�i>%B�L����u'�܊Y���� p�����o~���E�'� �$���'0��'G��'Ԏ#��Y�?슔qQ�ۭ0��z�'��\���ٴD�8���?����򩆳vwHQ"6�ޔ.��i�$�ԩ[���!����Oj�4��?E��	��^��2��L�"dq�Bфy� ��ԂFs�Z��|��	�OB��I>A`J�,�N��S��=�+e*ݝ�?���?)��?�|j+OrXn=��Q2���q����P-J� ��0±��џ�I��Ms�bǣ>a��`��$�/ޒS#f�Q�ā�P�����?�����M�O|��d��"H?�ɓӫ[4�q9�J�~˘\�H`���'��{"�3R��(d��:��Mj�a"uC�7���6�f���O&�$.��MϻT@m��X+=4�xu�X-�FhK���?�K>�|ҶL�M�'�f��C	�	�,<{�C�"�P�'1�� ��r?�J>/O���O��rtm�@�0�0�!X�tR����O@�D�O��Ġ<�$�iJ0l� �'2�'��E��$9�e+�O�x���Q��y}B�'���|BBǟe���k�&�H(�f
S���DM>l��n�A:1�F���D:J���6R�~l�UḩD#Vu˄���v�����O���ON��,ڧ�?�$S>0���S��tS4����?� �i�2�(@�'�o�>��#�怛vOY6P��P�i�sf�	ȟd�I���e�঩�'�,����?e�C��*(���B,�L�Z# #�}#�/^���0��O�O-L�r��2ӺeK��	 �@�!Ǚ4���0��=F��	U�˶
�~a��!w/XI8 #C�j�d��#o�\w`a��CӉV�(g���*���R/kRˁ�ND2������7$�a��H�k�����*�%��#���
B�^ev��b^�2���J�w�xDK�ǚ�� �#�㕢>)��"� �>AT��b�!W��KӃO+,��T���8ʰ��1枴*�DbC"�4]9$y*�o�E�X�f�6D�.�RB�^�U�zU��iE�Q��[�Β����Iğ����?5�'����#!K�]kǤJye��8��t�B�D�O�[�N,�)��:%n�8��(a����|7͊0<��d�O
���O���<���?�� �4S㏐$a�6x��n)?b�w�i8r�x��'�ɧ������t9n [W�׻C�SW#��8��=l�ş������uy��'��'��� G2�SCS�� 	Y/�O��#b�+���O����OR�`D�5r�9$eZ�h�}��%�Ħ��I�\ݦ��'��'0�|Zc4�����1g�]�&�N�vb�p�Oh��F�:���O$�d�O`�r��QJ�H���5��m=���Q%���O����OT�O����OX]Zd� <ڪ�3� ڰZO�� ����LX�O����Oh���<�7Γ�V�Ǖ7��)��	�rQ�X�F���4���O��O����O��g/�OX�����aĀt��)�1S���"�	y}�'��'N�	/�8	�OJ�L�)���qe0U&�UC�e�]�7�O�O��$�OnU@�+$�	9OR�X�
�? b%)6b�::bf7��O��$�<��ק���OL�D���8��.BD���E�(P���P�P�����		g�Y�?�Ol0x (U��2�
w/����ٴ��䑈V 0���O���O�i�<�13o�HA¥�k#�C�+�'{���lZߟ��I(i�^�	o�)��mBƬ���Y1E<x����7Q�6M�8��d�O���O��ɮ<A��?�3��A�u�tEο57qCDJ$]:�V��2V��O>)��.x��q��	�!�V!����<��޴�?A���?A�ȧ���O��$�O^���"LE���U79ܵi��ԖW��c�!u`Ta�I,���0u����5�Wn.��:�툧�M�|`R�+O6���O��D(����l�G��6V�+�)Lr�Z�p���RH�	��	ğ��'�H�ӆA);~J� 5��``PU��a�?N�ş��	矸%���I矈�sZ�?����lK�0B4D��M�����Iy��'��''�	�%p��Y�@ �g�E�+�Μ��>���oZɟ������&�������R�T?���T�����V�V᪬�e��x}R�'���'�	XSrp�L|��E 6CنT�wkߕL�Z= �W�0{�f�'��'`�i>���j�)ݓx!��&+vS��ʃ�$t���'���؟d�g�	|�d�'d���5��%ې��Y�(�����)���?1.O��"q�i��&��%��<�f@��=@�`�	~���:x���7�i���'�?!�' ��7]�iblF�q�&�C�\�7��O����O���w�s���M�EX�%$���1@^�h�.h�%IݦI�G�����Iß ���?����iX�|��qi�!U�Z�2g���uSL��'V� {���S9.ՈT�RK��~@r��$̘�[RD�ڴ�?!��?�ף���?ݦOV�kU���(�0A�_(!��)��A�'Z�b?�	[?!����v�̥�&��,;� �N�ɦ5���q�F��'L���'l�z�fא\�}�C��d�,hÒ�#�dI�K61O����<A�1��G�Z�B��v���ԡ��U����OF��*��ȟP�:^��NI	Ge����Aߌ�o�}/.��?��?Y*O�k�͕�|�ֱe���ì֞DN�t��(Jy}b�'��'P��џԗO���,>EsW/Ù_Q���Ț\����?����ONMB�K�|
���ML�i���`��x��!��:������O��x���&���aIZ�i�*M�P0h�q�mӜ�D�<����
��(�`���O.����|���+R4��e'�4�&��5�x��'i�	�h3�#<��Q�T�	$bO��@�C.�;D�H n�Jy"-S�r��7b���'��d�=?9ad�9v��QM��tp���ej���'�'bN�~(Or��u&'R/w>=���n��sçj�Dl�4��O �d�O��D柎�S�4'҈J���`e�N	���h,I=�v��L�Gx����'����5��+d��I�W�[ Z�H�h�f�b�d�O����?���$��S����	B3ܥp��P�P	��'	���|i�4�?a����$NK��T>9�IM?i���>�<C��yLHL���ݦ����&Njؔ'��ꧧ�'e�H�%W;���#I�)f�Du1��,�M,3��ڟ$�	ȟL�'�`H$P�@��P�ɇne��j�J�D�O��d�O0���<9����HV��k!̋�o���7����MC������Od�d�O�˓/hp��9����ƥ ���?3jzrX��I쟐��Sy2�'���؟(�4o��B=3��t	�"E��h�@��'�2�'f�'3bl�Sk�7m�OR�dG�a�,�3c��d�,@@����٦��	����Wyb�'](�НO]��O�Ag�E Xn�qz0�ђpr��׻i�2�'�'�
# j6-�O��O^�	��3�1��$���F�Xo�㟠�'7�#N&���|��M�t���&�S	+vI��E��������f����M����?��R�'�?&ʢF_zE�#��S��<aj�.V���ߟ���MI˟��	cy�O-�z�f��89���iF�[�[:�	n� 3Mr��4�?���?Q�'�����?���E�l�gg]${��Y\N8 ��i�x�zv�' �[���}��d��&�*pBv�`���+G:�q��7�M{��?Q���:q�i���'��'7Zw �%���2Ir@i���P��н��4����O���;O��ȟ���ڟ �V�Eӈ��aC�%v!pDx��ש�M��&�άy�i�'|��'��'�~
� �Eg�[\La�Æ>q���IZ��ۅ�a����ҟh�	�� �OJ�Q5g�> #�V"o- �W�D.U{f�s����OD���Op�O'�I۟�
!K�8l]r$�B'Q�w9D���1:E��	by��'�bZ>��I��ܸ��4q��`�c9a���HC+ِ �1�i:��'sb�'1R\���I?�
��u��!J:��:c��H�6�Ql}�'���'��'�]��lӘ���O����O�3��$yGb�^�a�cݦu��ٟH�	_y��'�P�Ou��'y�0��A�2�����P��Dw�f���O��$�O���%�æA�IПd�I�?``g׌� U���t.lJ��"�M����D�O��Z�=����O���1�b��;^B�0ae\?U��U�{�����O��a���¦�����\���?��ȟdऀZ)|�w��+j�̉�G�
���d�O"ɐ3i�OВO�i<�dC��iC��"�_ p�C��M�eD�!PP���'r�'����O|��'^"k�I���3x��Xr��5��2�^���ޟ���O~��t�*'��	�@mP�.��e�.`��i���'2*����6-�O��d�O��D�O�Női
J�XZ�H����\����4�?I���?��<�O���'`"M��q0��Tb1!�*���ʟ2r�h7�O�x�4d�Ŧ���Ɵ��	˟,�����	24ȭhEϮ%Q��r\FC��E�Rx͓��$�Ob�d�OH�D�O �I։��[���0;�f�0L���l�������$�	�����<A�~Ҷ��Q� $��pfJ��h%E��<A(Ot�d�OL�$�O��d��*�DmZ�R��{���#)��r��)I���rݴ�?1���?����?!/O����g��i�e� �r-��n��cFQ!Ǡ�nZ��������I���)	�n ��n��h��¦�;��4/�Pc�,��wa>}8��i���'�Q���I2,��Sş�8���߬vS83ri�G
H�nZ̟ �Iǟ��I�[r��ݴ�?���?��'
��@��AP=̕�eZT;h4��i�RX����;|���S��p����45Q�Ir�l��n���Efϵ@�m��(�I�V�ʜ��4�?���?������� �ۗ�V6�NH�E>�@싷_���ɟ6VV��?�g�ɐfgb�r�ߝe�t��F�I1�6�
�p���oZ���IΟ����?a��ܟ��ɗX�T	@択Z$�)�넫?B-�۴U@������?a-O�i/�)�O�������ׂ7L�����������x�B�O˓�?��'�&\9�o�"!ԴY[嘣"\��ݴ�?Y,O�l�d1O�������ݟX9�eԢB�^�!��$>����s(^��MS��t���Z�W���'��W���i��)w�݉8(�]� Ӧ\ ��>1��Y�<���?q��?�����w���Å>b����Eܓ�����N�_}�]�h�Iny��'���'��[Q�
ef8�˓h�!o�u`�)�yr�'�b�'�2W>��&L��O;`�0�D;
"���R�`a�-�ڴ���O���?a��?1 �<Ia��M�ʸ�r$/P�}���P�QR�I؟`�I蟈�'P���]��'�?�$�^�Q9V��=�Dض��jH�&�'����P��🠲Rh�H�O�r�%�̄OJ�M��J�N��[��d�H���O�˓���RsV?��ӟ��$2��y�c�@*0��г0 Q�rn-دOP���O����>��5��?��W.�(jq�D�& �hpv�p���=g��p�i!��'~"�O�h�Ӻ+��-I#�uIT|���A�Eæ��I���z�Fq���	]y��)_�=�2��'��M�S$�+��H&A��6M�O�$�OB�	_}�X� ���d
0�:Q%K<$H�XK1�ɦ�M����<���?�����O��ٍh��!�͞ L�"���	�<�,7��O��$�O����AEe�០��N?Yv'�.@�A�
 rz `��OȦa&�܁�iϟ�ħ�?Q�����ۊ(�v�C�+_�$�p��>�Mk�7��롔x��'GҒ|Zc{�Q���%�l�[��I-	GP���O��r�?On��?Y��?�-On($e��~�pà�ۚ'���b�X8dS��%�����,'�����\C�!H#>[�t �,�̨��H*i\40��Fyb�'��'�� EF���O�)��5L2��z�h�r�܈!�O����Oh�O����O�]ʀg�OPy���2h9B�����#C��eCM}B�'���'Y�I$-�04aL|����Eq��PE�Z5���v�@3)���'��'S��'f�I��'�链u��ݣ4�*h��T
ܹ��i�2�'A�
/�LL�K|r��Z��'�4�Ճڢ�J@�W�ZW��'.��'��M9��'�ɧ�)�,�"Ւ�`�c��p���#���S�D�u)��M�X?��I�?y��Oj���Aښ�b����S3�i�"�'U�<���)�>~b�0�	�T/J�u.̧�-�Y6m�Of�D�O��)@�	ğ�,߼�&A��	�A# ����MS`O�<�L>E�D�'�~���@�4�:��&M=_�T�ˣ)tӄ�$�Ol��TxĈ&�������d�����Y��p�%Q5��Lnt�(!�1�L|2���?��j���s�^� ���sC6q?����iHBX�A�hO���O<�Ok�V5^p��Bկ.�1E�("d���g��%�Iiy��'���'��	�+;8�������G��;�l0y��S�ē�?i�����?a��S$2/����r��q��Q�<�I��P�Iğ����]�|��	�42����]>+��qHX~ $�ش�?����?�J>����I�f,�� pa�ԥW�(y����`�)k�%c^���	���IXy�I7�.u�
§w�d�A+�?h��������	ݟ��?Q x�D�Ze���U���u@ە^�b5oZ������l�	�<�޽�IƟ��I��@�S�����r-�[�T��GA;��uN<i�����J(��ݍ�����L#���'�?^7M�<�rOE>~4�6�~z��"p����3�۸z���;$iC5|0HT�g����O��
6�IdܧMjDat�ˣ[�|���,���n��̘b�4�?y��?�'/��O�a�S��su�Ъ���V��`�b�צ�P��!��O��a�bX<P��,}�m�d	U+��6M�O����Ol@˷��U쓫?��'�2		�;H�	���n�Bds�}��B���'���'�r$ЋW��� �H�I�.4�q"A(F�v7-�O���"�E��?iH>��Nx~0S'D�"Z�ɲ�k�h��'�Јy��'��'j��?Z]���?=n�"��
\�������?���䓕?���i�$ �d��p �Ls$ʔ�>������}̓�?1��?	/Oz���G�|�nϑy����AK��r��@е�Dv��ȟ�%�|��ȟcEŨ>���B�a,` A��;w*8ȷ(�m}�'��'��	<<4�xO|���DM��Xc&ܼT7^�J@�4����'p�'h��'0j�
�}��!l�`s�D��*4h�M����?�-OXyp���H�S��0�%�a�5���м3���g�!�K<q���?��~�'K�IlzrmK��E�SS��k�?��]��X�ǂ�M�2Q?)���?̓�O���H�W�z�*T��'9=�ÿi���'�t�����7�px%,3�NdP bWћ���Q�7�O���O��)�p��L�*�C��֊A�ǷZ��"�^ئ��2*���O�"�3M������zj�Xr�w�6��O����O��<�*���������C�%�J�87m�=Wđ;3�T��OXd%>���ܟ��3N�*���JS�t���W�i��1��4�?Q��J>���'��'
R˧~�'�}�CC��E�l �Dퟠ[���N<�H>���?����?)��C¦-
B�<*��0GFcUҵQ M����D�O��d�O��O��D��芷o=	|�pF��utX�u���G�������ܔ'fRɍ��R�<����̅�^���W�z�6��O��$�O�O���<)������R���ޥ�ta�0(���FV�h��̟��IYy��O�p�η�a�O�Ɖb���15��5���զ���|�Iٟ�F}��W!EQi�i'8���Qˣ�M���?I*O�yҫ�K��H�S%��`�P�[JN��Ѧ̜���X�J<����?�O������l-RQ΃

�9H��={/��ʟ��E�Ꟑ��ğ����?��IiF�.x'��y&��X� ��j�ݦ���Vy�F 0�O�O�(R���3\��A��1u���ڴ�ݫW�i0R�'��O�O������|H@GY)r�J�
&�ܷl� ��	ҟ�� aUa=�qѧ�N�V��qπ�M3��?��}<��$�O$�I�!| I�m\,4h
��h̖t�6����OV��O@� %΃2[QR�!���l�¦a�I">"�K<���?IM>��O�2MC.iR�aa���4wmK�>�� F��?���?�.O��lT�S�t\pS�9:��1���V�P��H&� ����,%������)�F��������g�E�fi�a߀c��2��MZ�z�ˋ�)K�|0�������6�2�I�"�x�!��Tݐ�Y,o�PbC�=�qO�����E�L���h�7�B=��KR>&��DOF� 9 �#I]�����	�?u�T��4.�d0U�Kf�hL2��_vaмR"%Di�f 5�!9o�Ձׇ�./_xuaT� �A`��v�
�M~ b6�w�.����?`O �[�N<_ ��p�L�r���OG�z9N���'�*�:��&qs�aI]7D�V�r�'h2F�X��B��ɡ��s``&G
.��'��i��C�� 䃙�!T�8rѷ���I� a"�8!]��4�ϖu�N�!$���O�8+B�ӨV�iC2�T8;IܱKN�ʆD�O��D;ڧ�?����s���p�$��/���oA0��xB-�@|'Gܽ8~$I#��
�0<鉢)4X��(9t��� ��
W>!��O"�$�Ob���K9o����O�$�O�Ҭ8��5Ia�ИY���S�ɞ�2��U����
&t�1�	��29Jp�2�3�DP#��P+��)h������4��=0�	�,P20!�	�Io�* ��|bAE�[�fPg!O,D�(��2b��Hr�L:SE�O��O�X�F۹Q�`���$�ּCׄ"D�X)��S���Ѐ�8-�t�P҆;?yV�	���D�<1��2 ��G!3��EJ#�.e��p�Dϼ�?����?���2��O���n>���'�� ��H2`�C)8�ډ�!H�:���y�L=���hPax��p�jFB;�m���ǄP:�\���G�-���Q�aU���i6�\x��A��=5�t�b�E�*�92�E2���O��O���O��\���؀1*���"�ip���d?D�� ��"�K��!0p�.>��h��$�����ISyr�  �ꧫ?S�%t����D�u�R6�?����d����?��O$�670\�xc�>XZ$6�C(sd��s�ڿB%DţF�J�^��xr��,_��hv����=�c�i�hh���W9?��=�@�Έ<��\��������'��xK %�^ȧ霦�N�ٍy��'C�e���D�(g�x����`Fm!
�'�06�*x�i�e�msr���g/�ľ<9ӭ�!?���럜�O'L�xq�'���x��!@�|mC�c �k��3�'B�->S�����D4g�X41 ��O�SE�����F���"��O��EGZ�H�����&]�9�$�0�	O<�H�Rh���S�S��A�`�J1 ��r��>��Pݟ���F�O*"�	�)7*(�T
ߔ=}P�È���y��?v*�h��W38$AS!Ɲ�0<I��I{�ꭱ��I�Z���P�o̘zcB@��4�?����?��� p��3��?!���?ͻh��p6o��`��dBƀp�(=���]���J$�
u
@�QT,^��Od��'yL�$�.5�\ 2g�0e���p�ͼ>�����DKNGθOal�'�j=�p"ܠ?�R��!aT�tY��'9��>�^���'���'� bJ״e광�ʐ�A]�L�O�ţ�Ǎ�ְ��[r��񐜟P����?9�'�����F,<yU���K0|)!�M\�.�b$�'5"�'��aݹ�	ΟḨXq�\�C(�=MG�� ���K�� DV���ajw�W�P���-�(��B�J+�2����D(�Ĉa��X0$.K�,�1[G���	�%.bS�@� �|8)t�;��[�C�����ʟd��~y��'4�OHU�`��0�����ơ#/Ą�u"O�4r
^Bp�/g2ч�d�Цa��qy��X$0i�6M�O���-o��Z>i��j� �ku~�$�O�Z��O���{>MZr̟�U+lX'�<�$�:P��B��3XI����*O���d�[���O�RG��=�Ay3&�e��13T�'9�X���?���?a �ң[��m�uZ<��Ё��d�O��"|��GքpDl�`gᕅ/�H�7n^J<IR�iܶ|��E��+Ŷ�㇎XhHZ��'��7��h���|r����	���R�U�^�����q�Y"Q���w��'�<�D�>k��Egm}*�ʧIn$0l��(a��N8bx�O8�c++pX$��U�OVX=����� F�*�b]#1v��M���U��O��,�'�?YbK'8�1�@#$�H�r"N�p�<r%\'����J#{$Ip��c��
���
�6-bd(�G���J���O�@,�IMx��SW�P��w�[�����h/D���i�,cM��A��i�e�,D�#$\�=���1���9Â��X�B�Ɋ9Q���_���}��3&��B�I3=��4Pɛ�yy��o�eO�,�ȓ;��L*�J�)R� ���ŉ��Ą�-ɤk�+!`�U��{�6 �ȓ1�v�b!]�.$RLYo�>O쌇� )��A`��c���bl��V:(U�ȓ~E�H���)C�QB-�C):���V����IjD�hP̈́!t�@���	ۈ���NG,0�]�T�D6�Z�ȓ���S_$WT6���'[�v����ȓjL�R!�	�!r"M�6�C�	�+�Q������!w���0�0C�I�=l��R�òM۸l��t��B�I 
>��Q�c|`�D��?��B�	>8���@�'@m2yK�cC�4B�I�l��@�GT�n^a�v�n �C�3cĶY87�t�k�Jۮe��C�	 }d��:f�K3u?�����J�C�I%D$���7��	Me��Y� ��S�zC�I�I�Q���;i (D��n"'�C�I'R��u��J�[.����J
;��C䉂V�]
��K��t�3�U��vC�w��3t!��8l�]��@T*rmfC䉓&�
L!�,ʂ&��!M�p(C�ɉgxu ��qv~-� d�k��B��|	� ��w%P�N�@�#�F:e��%:����",3e�CVX�t�䈁gŰ�s�(�0D�Q�sO.O�9)�%�����"v��;�up�Ш@��� i�GdZ�G�Ǯh
 ��'"H�(t��	�-ٿ cL�0)PR�6�>��f���2�w"8q0��3�9�҉&-]�`��n��Dr�C)L�����RwFx(��*;K�'��U�P��ꋫ,J��+�-�T%SDY�<~�����Oƽb|F|b+#\P��g��[��ȺSK�`?���	)6!##����|:�f�[y���*�A�L�n��qF��-�(O���Q��f���o<f�*P!P4O�8�g�/y�aB�5BŊ���DA<挳��-,���,�$+�(�i�[������'�ȑItm�|~=I�oؠ{Zt㄁�W�@H��K�2�t��3�-�B�)#�Z���v� ڸu
���VF������Q�=�q�)<O������`�<�u�Y�P͞�r��^�R�J��<_�|���+�a�\��Q"E�T���!�:����(QN����	U���դFϊ�O���ńO���J�IPd�u�d�	iK�T�T���b� }ALRq,1O |EDB-1�����lX��J�)��C�eMF�I��c������<5X�l��4`�!)4�\��p=i��O�`�pX Q�Q�|vD�e���f�����%P��#iWTx��)��?�>}jVѪPE*�C��r�<���)=��S!�B_�+	JDx��Q%�R&R��)Z�J�.x���ǺD�*-q6
dC��׭�]��8 �asp��R��?���D!:f�U��:�6؄�*�
<z=6ڀ���R��e�Hm�qO ,�EAՀ	O��G#�Ș��WMmɚ�Ң�T����>!�1OBtB��NH��PCq,�8>��+-TtH��TG"��דN�T��1GA Af)�Gǆ�%X�,��FE�]��r���86��8����`NNY��%��:h� ��!P��E(�;� h�V
�!�$���ST i�R	�a<$�&(zH�H�Qg���NӠLF|B��A~�k7�܂=�|��a
��y�,��j&<	���J��3�T��qY�c��X��$��Jݤg���>)A燠@h��(",�(�)Y�<��P���� V�®B��+E�7�V��&M�*=�i�S�_DzpX�Ai��iRd�Ї�f8���!��D�^Je�W�A+����,�Y�YC���˟��'��.��|�)��E�?,�-D��#�a~Z����(~"ɰ2 Q6)JJ[ ��^�F�J>Y�����ڠY�)+ad�c4z<A�ۢ����QhĚ ���W���#�0�(��6�YF�hJ=?5��:6S��M3�M
Fx(P��|G�U���1�Ȉ��'N��9����hf0��A�i�Fy*T�<"���H�;b�*����x��c�!�3Խ!���z���o��|:N<�@)πr�IJbj��@W��2���/�,B3�&��h�f�	wj_�
6����k�/=��탆o��t���'�����(xv�K�bN�6����c�}���2c�a�����3f��������/��9b (U�7K�K��܇���:�Ƙs�J�pg%��JH}��皎s1l��kQ%SD�3�3?���&T�>���2t
�XSL@k���i��P�6���'g�q��б1��T��1pƥK8�H��-{<�K�N1Cg`]��5.�xxV�_�WN�(!"�\O+��cB��#���{��2b�6mD���酣_�I)�èb!Թ��AJ�,���X -уJ�Bᙇ�ݍ-�!�DE�Nv´���FGF��V���`PTŪ�/M�~�l jpl�
LEʙA]���+��OF��R��� �TĨ��&?�A@�IS��6r��A��z�k��I�CEl@2\����O�Kh�@�C�)Z����$jp��3�WP���I�X�P���D�a<r������2G��SK[�B��6�2Q�qO�m��C��Q�>�;f��Z�ER&�Ζm�����CC��G/< �qŢ]5t#2i�4h�P������*��TA3�'� $S�.�6_gf� �S�&�A�'A0d�l�qn֌A�<d*�i�=B�����7g�8/�Y�i�@ITM���7�LQb �l�Z��ֆ���xr���5�^IX�c�=���˓��O�Yᕆq�f�qO��ɾl0s�،QNhsk�}?��ɗ��6S����[�N��p��a�	x~>�����̰=y���S�r1l/	:HQ��4P�R���o�"��eΊlBg*��~P�$)�>I�HS��fB�S\w�<H�O&�*�����9���@%�`#��'�.� �d�o��
�i����WͶu "	\7^Ruc�CO�@�D��`C7@R@4r�-E����?�� ���~�µ?��ŢeR1Mf���dȁ��'�880$%�M3�"'XH1%��q�'HW����͉>��7��&�F+h��\��OM3#6�GY	�fnC#K���9�(	ֹ1m��+�f�Y/2A#m�*N2��̦|0�Ok��k>������L��yQ凨z��a�b��m���r^��1>��O�u�=!�iY����҂\���Q�Z3�݂FƼ�شOdؒ� M��~b�v����l�iqx��B^��=�%�!+�L�o�=z�X�{$�n<0%KE��y�⎖�'�P3b��s�2��+�h�z&�i��{fF�.J
����ͭ?� �5�%�R�J8e��2O��x�u��C�o�p�[S�iVRS�%��0Dx�s��{c��Ɉ- 2��������3Ɍ>�?&K�<� ���;�鑳��MFxRi��YZ9 �g��D�\�4"�?VȘ�t�z-�D��K]�E�E�����pD��2��4*�?F6��q 
�۵4����յ.gxJ@�`�\I�F%�I��4��� @�c�L@�E��r��H��J
/� %:���>T�0(N#���~���XM\�4�c �&2��	FHN:I��	�XȅC,	}����4N��j��]�0�:q��ՠp�%�T�X$A�W�I�F�X%E��b�b@6[ 	fҟ� ��CFЍ(s�չ ڶ�┗��U�B�3��l��!_2�Mse�!�J]isR� �ʏ�)X�d�"|��� ������E�L �Ç,�H�ş������G�,�.𡓩��FdLe�d�8y|e�����u�Ӏ��,O�e�	���,Or��P[�V5\����Ør�T :�(�+NŰ�iQ�ջ�p=�;LP<�˃l޸	y^�tTU�|�	�TQ��<�ɇd�Xy��~b�P>udP�얈팠@����0<�$�7$7Djc�<x��` �Mv�	�dܱmK�a�%�"6�P� �lW�P��ٲ,����vݓODS�n jBp_��*�@���w�m���`~�藱ant������)6�E%��'E�lCD���H�V�D:�HQK��'��➤X�lB�g}�b�(�t�z�)W���@U�p�V��&B��r�����'��W%��a�nO%)���'ۋl'�7��8v�T`�J۠_��������y�WK�OW0�أ�HRO,��O>���,���E|��F�<�g?Qg-K s6b�˒�h�fȫ7,Z�'V�2c+��l�@ ��d��:C���'�r(q�G\�wi|�+�/ڨ0P�%�#�2'��O���ib��I�N!?QF���&�?*�e��(Qu�L�#4ځ
�c�PtH�2��E8F��0a:(���\�@�*r��aǎ=�a)^i�8�	�b�̭r�ȓ_"�n�?@�3.#\Q�2*��Z)|�0�Ԍ=�\��6�%m#������m��02ỉ���^�c`�J������0�f�_�L<�4;�	֋t:z��Ǔ?�2��;=u#� X&��Jl�u�O!:��^X6��H~:*�:��Ġˇ�4�U#�>�t�Z�.L�X">��	�&1j��㫌�+�D��!�<�3i׉i���;�f
&Rĩ�"mɬ}v��O��Q�Mʲ�:5��4gԍAŜ���\��杻���I�P����yRfΙ�x���N�2�L��(O�$&I#R�H1ɼuS�hA���W�5 Q�_���Y3-�64�8�xɟ�l�@l�_��鸠/� 9���G"��ND������n���tIO����'[
�1ƕG�=S�-]lu������0[c`]{@��S8�X���J�;��J\�����O#}"���(�p)�f�O���BR-JE���	ڿ;Vp�	5�M��az��=k�����.�&!�Q(�H,t|@�S�'�sq�ē���:1O�ő����B�5��Q:�?	���]�{Z��3kF���Y�rkŭO1O�X�vcՍ��$���(x3f�5�>�3��YH�kL#8^�E@����Xq27 �O�5��J$D(x�h�e>YJ��	�d@ai�/[�6<`t�'#O�Z�,�JR	�fz��h�V�>����S���0�ɞ����D� 0ԹAY!#��[���NՄ�,�K�T��p*�[oTL��	Ǽ��K��S7)V���*�Q��^��(XqN����v�*"B')șC3�/�7mF���E1Q�8H�D��1��il��`���;a�����k��">�d��]��qc#D��b�0�eE�<aK[J�DXr�S�6�&�j���k?Q/Ҳ#
�/�R��c�Z*)F{����[@�Â��������_;�y�l����4��;8X��q����ƈO\���j'@6����S��)Q��E�8+F�sl#�Of4�DCV��<(���r��]:�jV#�dT�t�'N�̻B-�h��`ʋll̫�b׆$����	;[s�ڱ)	|�
��mǉ�Z�c�EiZ�`*�ǚ����:��O+�,��%E[:�Y��n�|`��0���`��#g��5,��;�4۱�%v:� �%�(���\�b3��ӊ.�����0�4��_�B�	=1(N@h��
�z���'/�M�ĈY8h���4J�Cq��#pJϖ���c��#43O�>���g}b ��L�pÔ/sɐ�h�,Ǌ>b��P�F�L�0�	�&Kr��d^�IY�Ѫ3g�e�$�r!ŭq�t���~�6�[bW�ě�mS�r���ٌ�Ď��v a�狉
R섂$@W0�0=�w�U'm�R`P�#�86P�zRg�z��P��Љz�d=�N���pۤ��)E�
���@�Cy��d�+�������y VĐ����ZVP�3�9��'�Fq���a����jU,I�Z��}����<L�9j�Mԟdl�$�"��sy�	����Ě�fN6���+��(O�z�O3G���/ۨ��q ��@�#sd0qХ�q����4J���i�n��4Иq�������NT�6�Y�--���ΛmnD�kg�1�Or`C �R���H�#hE����i �A��BQ�s:ʓP�� ��*�?e���/�,H���N�"��$�܈�䅾wTx�z��D�J�x�Jq�����/4�*�yʟ
	*��}�Āx��i�x�J�v]�uq#a��UҘY�s��T�� p9�n�<|
�л��0|��T���@iv���H�{y� ��`^%�p<�NP	w.x	we
L	B�Cq�T�'J�q��X�k��aH��[��Y�4>N5��N��x��([�G�:Z����GO���F�W�C�"}�@�J�@��R���$E�Q��US�?�����T
O�]6�)8�`8D�8CaP�?
@��QJ@҂�^��9Ai�<����:YB-1H~�=����2|6��΢2�a�m�<٥i�6	r�	H�U�:ĺ5��O�<"�ؽ�ޔ:��B�I.���IHa�<��A�7�l%rAD"L}��˘Y�<�H�2zo�p��)ڈa�n��3'~�<YȌ�;�TA4�ۨv���B��w�<Q���&�������Qz�� Sp�<��@�6X��K`�p�sB�Wd�<�bS&�1�D�\4���')Lb�<!RנN��A�@ObPl�+
z�<i���Z?�1��Y}Z-���L�<� �J�c<V�x��C R9���q�<���Z#^f������AQ(�[!��m�<Q��av�$+ �>7�ml�<���v��%�D^�0U��� i�<�f�'�h"f�D���x�S��N�<y�O�;:���-Ѓo�R���c�<��h�� h�q�ѳR�а`^�<�g��� �����LqSpXc�<	6l]5D���t�̀}�n�"q`�T�<	�K0)���J�4(a��H�T�<�`!��w8n���e�W�>�i1 �u�<a�L��֨!���*���q�<YA�'5���A�SѲ`zӮ�b�<�E�C�qE|�c�E�����f�<)��R
f����8\A�ـs��`�<	��̞T��q�J�.[6�<��#]�<�%�N�dj"�H��i��#�EU�<�I�)T��� <:@&E^S�<�V��L܈� ќIi ����G�<q H�M�2qR!ͱ.C�� Be�A�<�tƊ�T<;q�,9��I8�JO~�<�ä�;Gڼ�G�V�?����e�<�ߣt� �疤S���b�<	�ɀ�>��a�J��V|�D�E�<�"Lĵ�8�E���M���� P�<Q�흟t�,�jUAѷm�D81�P�<�%�b֤	0�J@4i�|9GgN�<�2�]�C���Y&m�-����U~�<�FLU��`Á��p���K�c�}�<3
Ċ��d��$YJdm�d	�}�<a@��%��c`�?Ҫ(D+�}�<I`!S���V�<(�ؒ&�}�<�%���{����`��D88�[E��b�<�nYm�$��bDM�d�Q���H�<!0!�>�Ա�D�1x�"�����B�<��Q�5��a@ `J�6��E}�<��3	r��ֽ�!!e.��B�'D�X������0� �Q�
��p�!D� I7��  ��%��`8��ҧ+3D�0 &��;n�2�;Q&	�i���/2D�Pi�KH�7��4PK��8��$�,D�[qd:ci�c�Ɵ���ۡ'+D�� $�'ep��#�K[���r�6D����/�����!��$�Ȑ��3D��R� ��ޡ�U&��R|���o0D��c/�:u����3	��^[j���*.D�px�2"hR��UHg6���-D�� d�pwC��@��ЀG�e�X��"OV�ӑ��HY�岴f˩X�vM��"O�L�Ǫ
��-�2��d�b=j�"O���˓1�ؤ���X��8�"O��I�,�1(�RCA��|�8u"O�B�i�vf(}i�b� k�ހ�"O|cO�	�d1sCA�D�{�"O	U�_�Q��1��h6q�"O�|"DcQR�A[r)��%�] "O�ɩ����I�T��P����e�r"O� �
ΰP�����%Tc����"O�)g!J�6��0�d�#g�r���"O����C0����e�5��L��"O���H�E
�D��DI�	lf�0B"O\��q�ӱJ�VJr�_�[d���"O�u*�Sh5Z`ʰdμ\�>P�!"O�ţ�
�[�Vx�p�B�?�ƨZ�"Oq�©�aݚ��)�	"ʬ8��"O,1�խX��.�I窅�qP��q�"O��F"҈_�H5xp�6{M�x�"O~�0�ō�w��Ȼ�JR�a�\�!C"O�}�͔a?X٨�i��!�X���'�ў��e�Wm�� ���Ft1���>D��g���j���6$�@�%m>D�l V�a�(j6DU9%�@�Ҡ�;D��h�B:A��)G+<��
�O$D���C�>�zPJ�<���k&�.D�H!���|�x� �+�̨��*,D�z�͘v�ݣ�n���
��e5<O"#<i�A��!<̤y�h��j�80x�Ąn�<����� �� c�A�]u�)x����<T��q�ޭ�U���u7P��Df�<yG⛌=�V���T�V����@-�}�<��b�&M�.�����a�����v����'��Ԯ<CWB��n��1��'��ဠ�72��6JL134�h* �>i b2�S�'*I�	C1ѧ>�8�U
��L��ȓc5�y���V�d�X�TBJ�w�+,D�d�vG�Yϊ����a�8H�T�<D�\b�c�"np�	�O�#�8$�!-D��H�E�Oڨ���*6�+�(D��RQ�F7y�8D�a^7�*��v�8D�����1Ī�S�]�<�"��c�7D���6fN-�iѐD��U5D� �@�
&�*|R,�:v.���A&D�t�S�֦�,���#έR�4��B�&D��s�gP�\��}Y��+r�����!D���ƚL����C��[r- D�(�b�#w�t˓i��z���k'-=D�<��Fͨczųt�ݦE9`�b�<D��@�Z*����KDv|)d<D�d�'X�-O�ᚕHٟw �M;Q�:D��r��Y(/���!�;��Q#�3D���0#!e:x����j�X���+2D�X����@&j�!@+��)� �/.D�
�]�j��v�F>4���x��&D�|�r�T?-<<*1�P��(D��i$A˻�%JU{24�2P��DB!�ą�5�.pP7-��n���+��[!�Ą�	���@�ģ'��e��_ %!��0��B�N�\�B�C��!"!�J�.j}��ߌDm�Q$-��9�!��5q�ݹr�P��p)R��9c�!�D��7�e`�,���vD#�Q&s�!�� 4�����#��ж��*Ep�
�"O@H ����\�x�+�%x4q�"O*8�"�Ǉ	�d�#�"{�����"O��i��(X�HSME�O�~��"O��S�O� �:Q�@�(qAj=�u"O��Q7��1m�q�Bn�$0Ơbc"O(\���..���#��"@-�̊"OB��$��'k� [�k�?O"�pY�"OF��w��+����.*R!�"O�a2@�0uv����9
��"O0AH֯�51�t ��oAe�h�"Ob�J��ő�d���`�9Oފ��F"O|���S���1��=w��"O象f�R&���j�B�0]ʱȢ�'��O
D㠈�&F;@��H@$h�p��"O�W�K�	�L1fϺul6=[�"O�|��j��B��!h�L�Bm�P��"O&A1���P�S$��V�*$"O`�q@�F�d��)n(~��"O�pp�[�Xf @�L .`�FUD"O"���X���Q��쉥 �H8��"OV��U#�S���𗆅��d���"O��
�a�+J�Ҝ���*<�&�;f"O�7�T
�f=10D1��4"O<�{S��$""�m��
J��XT�i��d �dd&�F�D�5Ǥ��ă�b!�d��n@`&D�����դ֮IC!��Ó?X]����P�,�c�׀�!��������,u�h0aL'*2!���ƅ�Ԁ�O��h1٤
�!�$�% ��Ԣt8�h�c`@Za{���D&f�'J�����
d!�-#f!��ý4G�a�t��Cj`��f��AQ!򤍴,'a��Y��j��G�<!����x��U���{q��!���-!�d�-	2�9pUN���%پ-!�$Fe��`Rj:K�*ǟ�!�!&��}A�bZBG`@W�Q<�!�����Sdb� .�u��;�!�d�vi���+��0�9o!��חTK�@�1�Ǜ6n�
�( �W�!�ǒJ�6x�P��!8��JƇT'e{!��̚�ʆa@�	�r���"h!��)O�� (�
��)X�䕞Qf!�1���beC��I�A!`d\7V!��7a
!f�Ĕqנ�Q#v�!��q���7䁶+ɖ�Ap�[�i�!�d� "�y���0²@A��M#Y�!�!$@� xt$�2\9�"���+ !�$G���hI��P�h�����ؽ{!��~���r���jׄ��T>U�!�^�}��꧋�U��z�n. �!��d��u��P<�ҳ�Vk�!�$�)]��-l^�a4c�'	�v�"O�t�F	)6*:Ѓ�\L�P���"O����X4�䐗!N+s�$)�"O�q+V�I�tT�$��t�^�s"O|���YKI2횅c�I� ��"O��*������OކH<̽�"O�\��dІ.'TI�f �<*Ў���"O�<Z�l `������~���Z
�'z�X2s/�b���lD?d�|9`S"O�}a��I���"Γ�o�*$*��>����F@5p��ٵL��-�dHV��!�� vbqML:�� ���;p�%X�"O��ߗ�,u���ًIj�
s"OR��gM�aRQ8���?LԹU"O��ӣ��+W7� 2�`U�G�P�a"O��� ������Hz���"O�8ڃ�]��"-��Y�(\�aB�"O`�3�!���hU�^�^M�ʦ"OZ�i�m�Z�\Qw��"^L�A�"On �gf��w�Z��e��rH.݋�"O&�����U�\qj�K ;X;VIAb"O��fȦO�"�@�ЋP5�i� "O���b憆�P�[�"?E'騃"O�QD#<�����y��DA#"OxpТ X*u�nY+���Gbt�+4"Oօc5N�' e*�j���1c.V�iQ"O�h���E�SU�$;��
+=���z�"O�Pj'I�b�c�ùQ�fU"O�9%�6�|ٓO%�&0�"O(z��-qk2x�p��4�j��E"O~l�+�d\"O@�2��0"O24�ȅ@ɦPq�0�ԭ�S"O�=�$%m���I�� �xT��� �Py�KT6|��K� p=�ԋq�<q��ِ ����>d�����A�<�ȋ2=�(U����'�޴O�!�$ݸ$~{P�źY˼�3@��u�!��Q�2����9�J`��4%�!�d@�>u�ez!j��Ht���Vw!�ĀY�9���!8|!c*� q!�/�i�+Q>D�6A˰ɕ{�!�Ę����B 9Д@�7)]*!��;/�|E�uM	t�>��c(L%@_!�$j,�])3��92��$�aHC5(�!�Ć�A�`i���G!x��-�ǁ�w�!�$ �,b�y� fa�e�ӇRw!���-z�E��/�-bq2)�� 9!�d�1f�LI��	Gj�ړ,��[!��b�mA�0j �Z'bT8X)!�D��5+h�z��̴LW����!�dA4T�vu�Wm��C9�q�qᆛF�!�$�.u~XXR@49"��䆏�b�!�ϯe��Q U��F�@��&@�)�!�d� �`�q�ңx�*�@���2z!�D�_��h����rFcC.xG!�Зf����>>�Nq��� x+!�d]�#�x8DfX3H���A�"N�  !�䆋0$!���0�|��ƀQ.o!�k�f�W��:8��ŋ!�$M��X{�o.Z� ��B�^�!� � 58ǌ�5�D��*�6a�!�$�)������[⦩bã�l!�d����)%�rFHjD#W�P�!�Ē f1XL�4���vi±[�lI��!�$��,�v/F�j>��B��;V�!�d�+l0plB���:3�ٙ
��!�ќG������4J���h�&�!�_��*T0�bIs"�'�Y�!�$f��;�� /[	܃� X@�!��.���Y&��# W�8�&�]�!�$ãB4ؠ�#�7��ٰNU��!�ف� �ƋŪw7L�G��Q�!�$��N��a���9*n��eܸv�!��H�a$جzs	�2/�8ڇ#�q�!�^Hyh��"��y�=�!�
Ss!�� >E���(	ʄYg�WW̪�"OZ�h��.mA�����A�l���q"OF���ӭ1�Aj�#W:8�a"O��GN��0���kPɋ3 ���"O��{��ޒ4l�q�H�� �1"O⸩�@ɔ09����- u�d��'"Ob,����t�� �lM�S�6-��"O��w>7Xv԰�E���~���"Oe;W��"\�pTx6�4<�����"O���!��L|���c(�=�d@q�"O�<QU�҃F� ���
4j~��B"Ox��A&��d�d���]B�e��"O��Z�����D��mJ�h=��Pg"O!q�Ԉ�%�9(�\�"OĪ�+@�xS�E#�$E�lD��q"O�L����zv��Q�c��	'�"O�Q�hJX��0���&"�	`"O���B�T"WZ���a�^w��Y�"O�z)qh
ͻ��
k=��"O,|ɖnT�8p
հp��*oŨ�Q"Ol��ώ�*"D9�3�&��0"O�Q�`���=1�p"���'T���"O
�L�g�\)�A*�A���5"O:�3��ڂ.♘�I֨;��!�"O��O؅-0 x7	K�e�8�"O&L�u�İC�^� 5�@6(x|4��"OD�3D!ǬLr��FE�kaL�"O|9���7	�r9٦!�/Z���G"O�!&�M��rtrC�TIS�,��'u�t�0k@�+���sA�ώ-� �'Ud���O�C�(ɧfX+"J�X	�'ҚT�"C��?���
WkZ���(P
�'_�\7@�# R����m�	�'n�U2!ð{y �"3d�+=Jr���'랜��ɕLQ���qN�'8h����'�r�IJ�@fv� ���0&a)	�'�lr�oK�FJ����ۆ(�|���'�`�KAPc�y�I�<VG8(�'�fU[��K3��]��/N$SK,�Z�'6 �9����*�YrJ�Iqrak	�'ՠyxF�ƈ#}<��J�@�ݪ�'1�� �T BdgQ
�~Y0GPz�<��DB�YP���u��)FR�y�o]y�<��(�>3�hm���U���$�w�<�rbM7��0��a��1�R� r�<q�m͗c�Y�$Z��ԉ���o�<�T�Q&=v��db��t4R��@S�<�P �A����Ҋi���C��y�<!�T�p�A�ߥ-�r)c��t�<��BC3L:�%�"� ���� �t�<Q%��F��
��W
r��x��
�o�<9%�B�9h��ɽ�4� ���s�<�W�A���È;W�`I��X�<��OA2\���Z8"0V=�ǓI�<�"�GJ��ǌ�q@�0�BF�<!whɈX��1�g	(K9\P�7��@�<���x�QD�4p~t���<��46�B)� E��n��@�Zz�<�c��"Y���NG1C��C�y�<A���%�̝���+8>�{t�t�<)��Y w��`���#*	D0E)�Y�<9�6#��=���z�1��́U�<�3��!��HA�Y V�&EU�<�&�S�?[b��K��j%q�`$�Y�<� �u���c`Y���S�+�xh��"O 0D�Q9�8�PAN�+$`�5"O:-+2��y��D��/\3Qb��Ia"O^�kiPX�`�H�m�[�� �"OR�9�� �.4��Q�U l�\��"O���f�2BތmBwJ��T���P"O4hY�$ZI��9����Z��c"O��%AO�V��B�'�u�!�0"O L� ��v�H�e��?oV\p"O�T�be��8��@�(�r�\V"O���*Z=9�B��0-���t!�"Oh��-�/2�R���+ހ!٠���"O\ygKܠ6��@�6~�X��G"O�aP�F<L��v
^�J�d�ze"O -(�͆�.��P��>b��!��"O8�y��#bl�٢�ɍ){\�;6"ON�CA��!���'�@f�	{�"O�s��'�<����И|J��b�"O�,賯
3Qjd�Su�ވ;<���p"O|���LI��
�!3d��3����"O���A	(C�B����X� �d"OJ-(Ј��:�@���\�x�"O착��S�q���@ѪԈ]��Ͳ0"O�͹��<�<೰i� <z,B�"O���2$�26�8��c	��,�i�"O��@Þ.;�����H�ej�q"OZ�����E6 ;C�"U})"Ofh���QZT�C4LM���a"O����#U�_�%�/�:]P�m��"O�X�$�܈J�B�H0� ?�zR"O` jvBļPYT��3�ȧVje�"ON��s�O�&��Go+U��#F"Oh	�pb_EK���TCp �g"OVD�Ơ�LH�b�"ڞx4ļ��"OL�!Y_��Q���]f�a&"O:E���PT�̬ҵ"U�}�n=Q�"O���5h�nX��C+~�ԃ5"OX�'Ȋ��d(CK�^�*"O�2��[�l�yd-Q�)!&"O�<����2a"@3TL�/h� Y�"O��QS
�9_�l0R5����}if"OX��
1�9��a�2� ���"O"]�e��9N�̪"@�P�r�"O���J)U29��NV�&��{�"O��1�Ƈ�3�P5��NT����I�"Or�1"���mh���mW�7W][�"O�Բ5�_.f-ĩ�V��#�l�"O���&�t� �$\���mc"O0�:����r싓�T.hZ<[S"O�L��Bj�ذ�	@`p���"O�eS�a��7֬I ���Tb�X�"OH�s'�<T��{�I6\�'"O�h��HT��l`�F�[+(�[p"O��[M�s�P�[tŝ
S%��ZR"O��0l��`$DLu��i�y��"OR	���L��ՒUIU�\�$z�"O�ģ�EWB�*���M�!;U�u"O���̊�y���w�1:�� :�"O��%��d0Qs�Ѱ!�6x!B"OВu�� YPA �9v��Q� "O����E 9Q�lE���	�"�,!�"O�, Q&�\�P(Y�#$D!�"O�<��KK&)�4h��FZ��ڂ"O�Л��2q���E�͘g��Z�"O� �,y�� 7�����x����"O�	w��i%(9�!@M��l�5"O6�{�f��I�:��E.D6�(��"OF|��\E���i*��H�"O�1�7e�o*���v�6�P�'"O�j��IF� ��F^?PY�%"O�@r'��A�䓶�E�% t0��"O������,����#]�G����"O�l����%T#���D��?6�D��"O��j��u�<��[	���4"O�`���Nn&|��+�6f�D=b�"O��� �҉�0���s�fՒv"O�1������Y��K�+5��e�"O���G>�(�Ԍ]���"O&X� �:[�*�	%e�p��dS"O�h�Q�H-hd�h�����Y�"O8��	t����@�m��""Oz��1�;{Q��ڂo֒}�2"O�ӉA��`L�Q/K�W�����"O�q�a��1}ʮ�歙dsb(�U"OH��%TTđf�I�AoZQ�E"O��"W�ì[=��D0$Q�}#�"O�xt��p,(P0𥋑A4���"Oh�)�-�n�d(c�ϩZ(�$"Oh��L�<Z�1�b��B�d�r�"O��
�bL%ix6k ��
at�u"O`q"&*��"hp���#'�(�B"OB� ��u���a�t�xuY�"O<�3����E�މx6!�-�$�؂"OM	��ǟ��$�`&H,āj"OR�+�FC%eK�˗%�V��mx�"O��[7+�?Js"tBe�ppB"Obh��#ِSmd�:d�#ilL��"OȠ@ȜH��Y�U��YO1ʇ"O�Xf�V�J:,�VI�Yo�K�"O��RA��P��R#�AmN,
W"On��Q�VP4�. L(�B3"O�pp��%h�A�6� K�S"O嘣�Xt�\A��Ϝ�p��(q�"O�U��	��q�,����r�@	$"O���$��L�y��-TP>���"On�!��*Z� d���Qm4���"O訲���ZMf)KpM�++>})1"Onu��`X=�������(D�`"O��*"��dԸ�x�Ț��\�Q!"O2  &�.a����'�#as�Y"O��.R�a�4PӦ�{� �s�"O��ra�Xc��K���3����1"On@��"����" @�L+�"Op��w �6w-�!B��g�<�"O��j���x�= O��
�J�')��7͔ѐ	Bw����|�I�'|���Ƅ0c~X�C �wAح�	�'dD(p��)'��E���tz`��	�'5(Up�Ⱥ*� -��[��8�	�'����tA�h=Pԑ�۞P6�܃	�'�v}Q�FU%Sf�2rNș�'��s��D��&퐦@�bQ��'�ԋ��6,�-�U�pq�Q��'A�őV��;bP�@6��u����'�v=P&�'g82��Ϗs�֠	�'�\�b`�Km04�GG�6dЕ��')��d��,JV���Q떗 *�TY�'д�X)snI��F����� �)���W�j<
�j��l����"O��e��il�"B_�_��}Jf"Ot5����,�T� !K\�
����R"O�CB
�(eD�"B�'�n��"OP�3"%��6\�`��A��b�rY�@"O�åܑ�ȍb.B�dy�2"O(m�e�`C�ę�+�)X��x1b"O�I��
Χ? Z}��*ɳ.�V�h"OH���D��%� ����:v�d`T"O(|���7N��ᡰ-	>��q�6"O�q�G��v����A2��3�"Oh�����]�REiU/��V�z��"O���[��]�8����������MP:5�!kC���5a6� 5E����Tr���E�g;�P��ݵ6��q�ȓH�ά��M�*�J�!���Ї�_�HH�$�I"("P���j� 'i� �ȓ1b��@�@�x\Pl! E�/w쌅ȓ`�*�K��{z"�p��2EhBd��r3�P���� M�l4r�@-pn�I��)p�%x�Ë�.�(2��լ> 2�ȓOol��Eߐ{-N��p��t~��ȓ+�����i�BH2�#�6ˀ<��'$���#$� =r����KB���J
�'=��R����P����&n�l�x)
�'(0��6�@�d��� Ҹ~&R��	�'64���۝"����(ؠo�¡�
�'+.�Q暣f�mٔN�)lV��k	�'A�RD
�@X�#��>Z��$��'�z5� 늓OjBj#���J�@](�'�
MK4�
)>ܮ]�ᯓ$Z�XR�'�>�8���;{�ҹ�K�zX���'|�8Z�˺v�~�� m�(p7N���'�D�#�!X-t�&�"����V,ع�'(�u��N�:|��ٰD�{w�b�'����̙�`��eA
b4�$��'j�-IaT?*=aB��$]���S�':ē 兼�|Ph_`�x��'���Z�Dț����CWz6�z�'Ƒa�T�
�P�[�霣���	�'�� VՊ<��h"F�b���[	�'�Ѕ��WCکJ�gPS׈��	�'�b�9S��.H�V�?�J�`
�'���Ջ��b��#e�Ny��R�'�Z��ʹl����Tg�/��ر
�'Z(P'N���]���V#�ZX	�'[��S��*#��=���%
���9�'�f}����1X_b�q�ʭ{��s��d3�@�r�A3F�'��Xڃn�3E_0(�ȓvF�O��n�0��� �@��1��i[�L�$�$<h���9�ha�ȓNʰyAb�2��TX�W�\y�"O�y3C�%���ф`�.8�䥘""O2$+C��Kv3�P�i�:�7"O��r���-"�$�k�.{ �"Ov8)��O1Jɴ@3�kh��QB"OZ}�ޙ}��!�lX� J��h"O�	��DE�ƀ{E+,VĠU"O�������y3�i"	�"O�z���NX��3�.�C�"O�t���[�
s�B����l�h<@"O�P0�D�|�Bt�w&�bƮH�"O�8�@_�E(u0T��5��l�"O`\J�-GP�z!Ɵ6���$"O� 6�q����1��ρm��q "OH��M��x5�YI�����D�"O8���L
,����gֶv<M�"O�x�<�� !�J� ���r�"O�	a�A���Z�lՍd!��"O����I�rꐹ�D��I�B"O�L�5��~ۖ����d�� u"O8<"����\���s'��6����"Ob�wK��f��t9�� h�(8��"O��ه$Tf���X��A�.����"Od]�U���d����tkȪ!���"O���e�#P"�9з��:F"��Q��'6ў"~���S�>Y�Y ��IM�@�,�y�#�=+^rH�2H���Rힵ�y%��[�:�)�5F��9����y�-�=<���w�� l��б���y�bQ>�![�B�'h����!���yR��9g��5��a��-b�b�$�y"��D��1�Z2]8�-(1�G����hOq��� �Õ�] #+L�J�1�d"O8��`�W�n� i�
H�V����'�ɐ摖fBN�¤��
 Vd��'�0t��ŋ7B�~�:�b��zC���'dh�H9E��%:�$߸c9�]�'fb$��G�Π
��hZ���'�r)�))n��*c�>gs�TzM>Y����J�:T�� �(
	\�&�?K�!���<�ґR� � v�*��'�!�$J��=Y6�%ri�Y ��%k�!���SI`Q #3lM�(���\�f!���Jf�1�c��;WIޔZg��bu!���l!פ�9X�i�]�d!�$��*����p`�4"6�i�2���H!�$1Q/P�J��C
77 �` E�,,!�w�Ѹ��������2�5�@���&36%����|�Hġ�O\dP���{�L�Bʙ[Ӏ�GJ�i��ȓx�z�{f(L�nFr�{�S�I��Q��V��Z&b�k����P5g���w`�h���]�&�����a%��F{���H&�eڰfY�S�0��!]��y��������
L�l���a�8�yR%�*3�(��BN�D�L4�� ���y�Z4E��*��H>[��0��J��y2��l��)�%G8:*����>�yR�*y޴};����]g�Lȥ��=�y��֦S{���ǋ$BsJ��u���y��{�Xqe"�7N�x��
�y�@x���5�̌!�y�b�(e�D�q���T6� ��̈́�y.��`!Э�/S�D^�!Ə��yR�����鸠ל�0A����ybρPJz0K�/b���Mĩ�yR�̨d�<���&���U2��-�yB�X�Dz>�Bg�ϸ� �����yb�d�%b D��
8`MX�M��y"k�R��с� �Xy�C��yb�$-p@C���;l�83`�A��y�
B�+��qG�F:p�&��HH��y"Ⅱ#m���'�T�b��H�� ��y���-�R����,]t05�V)���y�Ļw�xT���]=8���(���yRl��c$�{�܉�"@`G�WP�<�D�=�>9������Pd�y�<� 8� �F]������s�p"O�(0�K$ّK�
�21��"OvE�4��}ur]��إ@�� 2�"O^a;cBHl���	#Z�eyz-��"O��
Ǭ�J����qn*�[�"O��s�&H���{w,S�t`��*O2�tEəD�A(I/!�<��'��<jEo�+n��y�i�}l��'T�ʖEE�@��R�9|��:�'ڒH��n��r�n�b	�.r�Y�'P�ⵉ�2�4|S�O��l�NQa�'� �2���/��h��ٗi�L	��'ENi	��o|2d�5��f��[
�'����0F�����»[�j�8
�'$�uB�Ɯ� ���h����'?&�B	ؙ%��6\#,Yy�'r�m[pcý@C�Q��Gj+Ȓ�' ,$*ro�7��B�N�0U��{�'�J0���;�x ӱP��1�'t.]��NK�(Ӫ����
�IG��	�'O:u@�ήDMj�pR�^1�mj
�'�t�@�W���H�F�*�tR�'/���(5���x�_�N�)�y�b	6���낁��>���� �yrc�}h��U�A�R׆]���ѓ�y���yB�����}��ѣ��U��y"mTE^�3�e�x�2 0�\��y�+њ)����j� �Zwk	�y��|���ʵ���޶0�Q��"�y��' =~��0O�?������1�y�oЅSNQX���k�Ĕ�@.�!�y�(
�jМ=�2$�>bn�@âm���y��G6E�����i�堵'�&�yb��)�����g6]�B ��+V�y�H�^=F�i��?Y�@ � L5�Py�#K)AY����lԨs�&H�w�r�<��]�>���FE�u����+j�<!WK\� صS6KA"$����Bm#T��z�IB�H�]:��.�vt(%�"D�t�7�R��#L�'
���� D�t*��ݦg��S��Ĥc�Jy�Ì>D����h^p��|8F!��P]�I�� D�Hy�@%Uiҹ{۫A�r�CDn<D�<ps�Ɠk��:T��X|� #8D��K�*H�#p$�=���� D�D
�e@�t�ƭ�@�ԕ)�,Pv�"D��1��ge޹R�c*	��1�>D��f#��^���kХqR�qa�>D������.и��1��,x�]�&E=D�Pg��*M��,����2�*�ѕ�8D��9$�n�Z١�-/�(��-6D����c��kg��s��Җr��r�>D�<$�Wx���������k�;D�X��Ư}BHDjF��U�써Q�-D�x
Cm��t��*��Y��,D����-��@_Z��'KFD2���(D�J$�F"!������"lG�谑�)D��Q�`��;t���F 0g�pC(D�̣�+�HiP�B9h��%D��w�I�[�`���[�V誀!&�"D�L;#E:4�Z����[I7R1�'�$D�h�֍N"�&I��$�:��0�'D��+f�k�Hd���� @Y6v�!�[p��qo�a��Uo
e�!�� �S��.(����*1x�"D�3"O2@YUΓ�<�,X���6%��eZ�"O�a��'+f�ּj�2u�����"O�����
*��t(��y�^T��"Oh�`fJ�3Vh�s�l�r�"OV�A���(9��C@�mzD�C�"O��F�S�r	�%���h;J�:""O|X�3g|輸	�K:탣"O����E:�`�   ��"O���a�y�I��ıU��� B"Of�Yc��Mx���?�p"O��2(�Ur ��)ѿoCN�[�"O�]���T�/.�ذ��Y���"O\AK��=;�J@[�)1��2�"O�hS���t2l(ReB�T�B�"OY���<} 	W��^��k�"O*!�.ɺW+n�F�Q� 0:�"O��1D Ѷ91��@J1�Xa "O�$����-[y�M����/�Z-p"O���P=)~���mP�U��0�f*O�|+��6�(M�ů��H9��S�'�t5 �4h�*`�� �t�<1��Y�"��Yx�Ǘ%U\���l�<��l�n�mSed]7a��$	4��_�<���qk�i���6<fMxq��@�<	3-�%zqb��!�4;��KB�F@�<����8��)#�S�m���3q�<���8>_v��w&�':�F��5��n�<�������@K�o�^u�.�m�<�-Y'ph,ÐӔ����-_g�<��԰ �ԡ��AJ9&���J$LIk�<��d��LZ�JFO�5Q��2���}�<F��Z�X�� ��^jY��
YA�<�A���~�p��v�K�>�<z'�x�<1�JUIfe�$��/J�4�ahp�<�+�>	U�W�>�&�ɣ��p�<��&S�B6��!"�!�.u� �@V�<!A��+
����Nj.�U��a~�<�ehCMJP����
,�f�� p�<��@^6]6�X�!��
� 0�"�s�<9b��s��H��Ӂ3����v�m�<����/��)G��(rDT|Y$c�<��E݋���&'�(��
`�<���"D=x1�d�B�:���;�a�F�<�@�A N�|�AGW94cfDpGG�X�<	v�Q0�\"#@�1r80�-�U�<��G�)�0�oE�1�tC���I�<	��+;���'O�	�6["gI�<�3�B�.��u��o�D��\�& �n�<�Ed�1Iې\��)��T(ڶj�q�<�&�W"}�w��EP�a)t�<I��:��xA ����q��l�<�S��N���r4��:4��q��g�<a�h@.+���f��$ �4SX�<�C� -�r�ca��qܲ`� NWy�<qC�G) 9�MZɛ�A8 {��x�<A�-� ր�b�0Z��9�!�l�<���Q�.��4j��'�v�a`�	k�<A�h�$t�s���#@*�k�Ui�<!C�A'F�L��T��)bb1Z��Y�<9�� ��dӇ���L�&�Q��OV�<�Rɟ�vR�C��%F.��u%Ql�<�'�W*!x@0��0B��ѼD4F	�ȓa3�$�Tb��� kg,Q5N�p��S�? ���ƈ�FF�U2����r�aA"O�5�'�˄�� %ռ��D��"O�q�!+_\�l9'�&|�j=6"O�����_�Y}����ڽN��Qc"O�tgR�N��xp��'�&�Y&"OT�w,��Q�b��rMڌ*f�"On�`C�S<����taJ�/0�(�"O��;V+��n����B�&74� ��"Oq2��I�ӖA�r��!R�9�"O��K��Z�3�a8��#�����"OV�EfAo� %��K�4J:j��F"OF��K�"�Z()d�07(r@�p"O���*�3S�F ��BN3Y.��"O&��2�3d�T��D�I�82"O,�����8�A�☭y��q�2"ON�:�`!2ar�ʎa��"O���E�s�`��EI�h��	r"O"����8�j�N V���"O�Tq��ј.$F������M��"O�a��T�V�T���]1%�qX�"Oz!Js#A�C �P���1dIb���"O�)�G|ႂ�+h�U���v!��9Vp�0F�
3�Z�y�%Ҕeo!򤆧h@����`ޜt5*��iρ.�!�D��]%�܉u�B��<�1�ݴTs!�DK�9�����Ɇ�f��Rg	�]k!��t�N,�7��/|���P��ES!��wj慣���`��4�(<R!�$L�s[�A�`�#w�d�c A��F!�$]%/���x�J*s�0qc@]�NE!�D��'C�tQ�[�x���U�\�VC!��+.�����=Ke<��a�,�!��"Xx�Y"G��6�b" ڬ=�!�d�k=���cF�h���ę?)�!���[F4����)�( *S)+�!�DL Pa�)�ɬ���i�&���!�DT�"|�ɛfh�8��kv�E��!�D&>7Ht�$�IK��)R�>�!�$��D8��B�Pw
��i2qn!���+����@)zO����� h!��%I�h,csA�=r>��Z�#��BW!�bzF�s�fU-a+�8Ă�<X!��ۆ_� � B٫d�d�3�G�3�!�䛦3��8�*+����&�3K�!�Ě�95y �!N?E(X��� ]g!�d�{�΄��ELH�Vd[d"|\!�$A�Jfk6�AB7�S��@�WH!�Q'�J��"��:	,DT���6�!�d��S
r͈���v)��b�
2+!򤇹Z�Z�'�6	p&��2!�$����B�R����T!��1s z�ht��
��(�S**D!�d`_<Y�K�kՂ<�3iݼ�!�dS�r�B4���ӎ_Ô���SQ�!��:?��Z�/])#�fp2��L�!�;�l�S1e�5K�L����d�!�;�^e�w��P'�1��T��!�DF)A�vl���8t&x�3&�^��!�ğ�j�t��r`��e�
�oګ�!��{�����h���Ȑэ��!�D�25�0�zd�Xx�P��m�;M�!�K.�ڴ�gʜ>	�ƀ�T��h�!򤛌A�dX2GT�l�⸺�F�6q!�$C=|��4:(A,i6~�J e>.d!�� �P��AO�	& }� �qE���b"Oa�)�/,��yá$��Q�4t�"O���T%��L�˗剞�	�v"O.mav���m��#�T�3�^X��"ON�"QDӤs�u�v�ީ+�b�R�"O��Q� C��0��sn@�t��ؑg"O�(+ޛ>�p��4��,�:�`�"Oȭ
���>�K1 ��{y@!�"O<���P+��b�ϫb_�8�"O*��G+ԥ?)2cGF@����"O>�5&V',Y ��مf�h)�"O��*��)���g��Jp�F"O�L����!`�j����3nJ��7"O���`�D]�V�Z��#�"OF�&�Ϋq)(0Jք�/W�\iq"O<�Ιx8�[N��=���u"Orp{%m݈j��!���0&�P[G"O��U�?k�<�����9�&��"O�X@�&JԨ ��@���ր��"O��qt�+c��`�E@�<7 ���"O�
c�D�F���1-G�l�}�s"OF�� �\�G2�{���[o�y�"O��s�@����[���Pe�	JU"O�-�W����J�QQJN<X�8�y��?c����ònɒ�''�y��^�'AJ �ԪTc��d�?�y2D�=si\p�����\����݈�y��ɜ0����O�SE�]��&)�y"�i1�H(N�"pRf��y�DJ2]օ[�A�GS�*�F�0�y�˘�V*�����9	R���Q���y�L��mHxl�#�&��$Y�)X�yBc mC����V�Ƶ�Ю�8�y2a��2t�ٗ`��Tf@a���y��>C�ݱ�,­O��b�B
�y���	=BFaK��InV��A���y�bD�`"�W~����ȃ�y��Z=9O�UѷdF4yC�B!�	�y2*M�Y�1*����m��,��9�yr�GC�6·�m��q9b�6�y҃�cC������>/��0`��Y�!�$F�^S��Zu�G..YL\�r"ֻI�!�b7 ��۱5'��O�l�!�D�� ����e\k��d!�@O!�Ȕ=p*В�Ī Đ$�-ʻ7!�d��8Ǣ]9?�XYa�.�!�ڤ\�q`�\tp���ש(�!�Ḓ$Ê���uaZ�r��_\!�%�=�OF�&��1���=!��Y����s�>[���K�F-!��A�bDҬ/��y���!�N�O3�����N<d*����ޔv!�F��aAHƫc�����	&!�$!{����fB�pb2���!�:qzu�0�D>S�͛�͊E�!�$��M������C����U� �w!��	` ��`�΍?��ĳ��3"!�d�9�4�G�� ���(�Q!��OX�ف7�H�vZ2�X���
�!��˟`F����
�ML��0c�_b�!�I�!���n��nQd��D.� OHC�	2Cj}��[�UD�H�g�2s\>C�I�"�R��ǚt:�ÄO_��C�	�[�`���h� od
t"A͞*!��C�)� �Eh�CD�H�▎D)�v��"O�ňV��!Y�V��p��-�v�Sr"O.(��$��d�άQ1��?u��u�"O��ڗ���t��5�p��4�╀�"O�DC�
�@>�[�+	b��`��"O�d� -/�:		4�:4���@#"O�:3훘J�̀z�A�{�XH�"O�,Z��?~���,$*rǕd�!�d�0P�N��q�K�`S�-�!��;G����V��ZE������!��}�h��G�/��):���!�\A���Ua�	)�DжLZ9�!��^�/ϊT�sh��ч���!�d�3=Ν10#ū�z%h���!�D dj�(���6��dѰ"�!�ѻI���p�="�Di�WK�B�!򄍨a�pI��V�@ P,�K�E�!�$3?-�҄�P�,�~8k�KQ)8�!�O'L;`H%�My.��@�0�!�dƧ3����^�
�T0�G��9!��Z$6���ҫºy���#���#�!�d&V'�Ii��ֹj��5�5�N�L!��YaZ�ߣ/�Kb�ۂB�!�d˱oF��e�("�@݀C,Y�Q�!�D�#��5c�%�BՈ���a��n�!�G[z4�g���f�8]*� Ȯ�!�Q�q;LI1�O�*Ռ��E)�!���}�n�R ύ�]`4q���z!�W�y��A�O��]�%�W!�D5w>���
��(�*�͌�G�!�$]��X�%g�24Z��6�!�A,r
ѓ٨!�se�	,�!�DӔL�ŋfM|z��1W� �!��I�v�	���Rc���Y�jN�E�!��
���'��(
��-�B��5�!�䁓hDPY�E����@#��
�!��[�J�Z�b��;�!���/���!�MM�8-�U!I�w{!��6���	�b��|:�K�9�!�A=]:�H�"Ω���c�L�=�!�$�Z�2��T�=��R���#k!򄉾	�0q��NP�R2���iáb_!���`�N�K��@���!X�h]� '!��Z,b�Hw�4b�`�cN��!򄟛_f]8�����h�{�웿�!��4(Ey)�i�(�� ��L��e�!��0L@��ݧ|�(iZa�[�!�$ĵVr������Y���JULV�!�0�^��JY�~(n��˜%(�!��Z-gW�x ��ƻn�;Dd^ /�!��8��=�b��>-�<"t#�� �!��V
 5`#Eн[!6z�OQAV!���a2�H�agO�7+[!�۔P���䌄%����@�R!�D��Ak���E�)�@c_���
�'�i�BG�����r@�,!��Y(�yb��ZbƬ�--�'���y�� ."^���jA�n��c��yr�הoB0U�P�#PS�\'�8�y��fP�S�� D^uAe�,�y��K�T���S-A�J�Lx�T��;�yR-�������;�dj���y"BJx��s�=��T#�`��y��� ���s
Ӟ;WНS����y
� ��
"`���<��:u��%A"O>���̍�t�r@/�!�2��"O�-q�"P�[�� $V�
��`"Ot�d�Q	X�TVlN!
��) "O�����P�,�L�#��{��}s�"O�0�B�kG��0���9l�a�"O�����&}����+-����"O^�(qI�j��!��j�4q�"�1"Ob1��i�13^�%)�+��D̂�"Oh��,N*CK����H�L�n���"OM�BoTF��a�j�?��Q��"O*������n�t�r�ɚuq�]�$"O�L@�*�$1E���q���h� �'"O�!�d��Y�@�(���7Y��X"Or�!N�l���☨"Z�H/�y���U��C�ѝdE"�h�"���y�j�ir�:#g�
�Z �;�y�/�BD"0��ɠ�7�y���`M�p�rl�=pए$�y�O�D�4�cs!�h�<���n@�y�l�,~0C�ʍaک�ʆ)�yҌZ�g��Aw�R
��x� Z.�y�*ۣ�R�"d�-4����Բ�y�cĽhR�T�0Z�d��7����yR��'��(�p��GF�T�vM��yM�Dk���	2�&�
�y�%"�*�@bOK�~v&IM��y��ˏ0��u�����{��䆒�yRi��U���"�{�2���bͧ�y�M$d��s힊s�P�Y�o���y����T$O��rp�=�
�y�K��8��YzB��lq�2T�Ψ�y�)�h��� �B{��\Ӡ��y"��)�1�rဵ}��(��N4�y���7F�����y�ԑ�v�	��y��!
nց��
3&�����Y�y���9N�T�RO��(AT9�ʐ�yB'��0_��=%���J�Ō��y��K$q�*�����	���s����y�*Ȯa�@-ӀΞ!{wΤ�0�̟�y�̚�^�$)��Lf��q '�L��y�JP*J�ݨ��W�SL�(&H��y2�,^7�l[�� N���[��y��T 
un5���Z�Q$X<+�����y��˿1z<���F�t��i��&F�y��N�����᭄�~���R�yB$�?3~`J�b
z�p,As�B&�y���ࠗ���kШP3T�ѹ�y���;x�n�[F��#�L�33�I	�yb�W%7R~�jA �1��\��-�y C�m�ļ�d�I(��B���<�y���|�p׊��''���yҥ�$�^͠��K[���B�X��y"◖a���ĬM6IQ�H�!���yb��
h��B�cV�TJ�$:m���y�⃓��ز�R?N�p:Ec�y�,R7�l)�G/4�:�6f���y�JQ F`=����<.�F�*"�y�h^9-�J�CB�ƴ#�%�d�ז�yBKX��Ef���}�d;�y�%˼TF� �vL�FA�Yx�'�:�yb,a�ڐ�N�/(�p[g��.�y2�Q
y~��PH�52|j���!J�yB䕘_.��%�0vZ	�֍�5�y
� B�x�V�f?Dq�DKN'T���G"Ox����Ւ(�L���ٔJD���$"O�u����#�����
O�	���3"O�E"��7Of����(I�r7
ձ"O�����Z"UC����q �]#�"O�P�7��5TevT��xa��j�"O<�02#�/V�<�+�DC�p��Ss"On(XD�ֳ{eX�Є$�Y��8�7"OBu��%��M���b�47�X��"Od�����1b�̒lH>3V.��"Op�rMI�;� @x5DӮZN�,��"O�u�D̉ dz�cp�Q�%<�D��"O4jA�	�=���sf�"]E(IQR"Ot�ؖ�:O�t���C�b�z�"O� �#U)A����^��xb�"O���Q�M�"Fb%���S�� �c�"OΨ��^�T�t0�e��y�ya�"ON���,<�L���<]�ĥ�%"Oh���C�d�$%��k�)K�:�Q"OT����[��,��j,�ɚ�"Ofic`X�O�\�;�N� ^+�"O�⋂('�4�̉'���"O�d��F̗�`����X*z�Q6"Oa!a�V7�H9�,��xL��"OH����i𶉸�L ���"O��[�$� ,������_D��"O��w7^�hKF�^����5"O@��RĈfˬ���k_9!� 0"O �0�G;5�h�$��0��q�"Op2#�އ�.qv)�>�fE�e"O�Y��!3�`]����7 ��A"ORD��M�2E::5���zgN�9�"Opш�
�e7y�0n8xĂ�b�"OHD�s�/4C`͟�Q��9�r"O�%Y�[�^�qpI�o��)j6"O>�z�B�-sV(����az���"O�����8��Y ��C�1yZk�"O��ꢡ�	|��ʂ'�z�!�"OD�bT��es4pꔠ�Fv���#"O� �3�D#a�츱��'�*H""O�d)�^"=� �9R$���Az�"On���(�1@
��dJgu��;P"O4ɢv�W1~)�m ���B�֝��"O�t;QIB�<�:D*֎T�+�X`٥"O��ŅmŜ:Q,�fw��1!"OlTy�"+"� Su��'F���"O���rN�(T��X씘j��"O8���"d�j�+I6%��<t"O8����Ow���b
A)�� ٢"ON��� �-b�4�G�-z���Su"O����_C��(��F˵F���r7"O  JgLΗ؊�c$,�N��h�@"O$�KR�W�D�i�

�eu|@�"O�I2&҇�`�Q�ɀgJ���"O(��dˡH��Uj�n�S����"O�]���Y�Lű�m�O����7"O�9*�N"����,��	�JI�$"Oj���M�= ��[Ť�4;d�3"O���1 T.I��i@cmT�`��a!a"O�u�S�$�Z8P��ۂ`�, v"O�)p��x���e3=h�e��"O��g��+�8I�T�Y�F��-YA"O�A���!N�4J͓$���� "O.��O6"Y:Ao�uP��`6"O�  U�f(��cr�
d\$'T���"O*�yu��M��QkS��W�0@bP"Oʽ�!�:��9BL��13f"O>��A�"����K���q�"OJ���o��u�����81�(b�"Oh-	5c�0\x�i6��ot�r"OP����ϵ_2	s‘~���"O�<�wꝂR)6#���d�E�c"O�;�%�"���*IF^r��V"O�,(���F��U�䈶"O�� ��@_���Ɓ��}OXP�"O�e�7�P3o|1p��W�s5��"OU��"C�LJ�ٱ���r���a�"O�ez��-,8� �ʭZ��Y��"OB�)�V-4��}j����B`c"O�$�FA�9N�
X�Caӿ9�3 "O�A����)I��h��β����"O��Y��LY(�`a
��|��	�2"OޘP�K��*��HS8��(D"O�U�P������Ib�V'��S�"Oؠ ��F�`��QE� �ԙv"O�=SVlH����@@.�u��e"OJZd\.��5
��Z�Z<�"O$q�q�\^�d��g�I����"O�H:�	��~��� �d���i�"O��`rn����@2`)3[rBS"O�|���Yq��0��W0|I�q�"OZ��'@:Xnb�`�n JHx0"�"O���d� )	�����	(B�V"O��SM��vT(���Н�"OҹaS��
Q�q�BjN	�y�"O�N
psZ�"bI .bdHy�:Od�=E��I�3+�d�`��C�)iңB��HOޢ=�O&���c��
JH��2�
�f�,!�Ox���Ҫ�<�Y�E�f����
���3�)�Sn�D�Z
j��f�3${�=Y��ޞI�!��I�T�h�#aLM�
��Q%*�r��d��0?!��J=P*fйCmՠ����B�h8�('�H�����	�F��#;��-�g�,D�,��β`Ҙ�r��Z/3�}@�O6��[���SP�h���K�:n�M����8DC�Ɇ)���4M�	/�8;�،O]4���ئ�K���Ӻ�$ʞ2���gl�*52���j�<Ypb��PrH�����"����b~��)§��e�@e�/
D,��Q�]�iX� �O>i!.��
ٹ��÷hO�0j7�D)|O^�Y��	9ҕ8��N�vG`�a��	t���)����k�iM <�0ͪ��0 �1O������֔P��[ՄܸDd��!�$�O���g��4�[T��i��ո"O�P���%]��%l�Fà�jQ�|�)��S'T	���6^���IփLu���D&GB��``	��2��S�-X�ح�'U�r��8
�G.Cd�(5E�6i�p�Сk6�O�ိO$	A� �������j=��q"OԄ�wB^�s�<�.��)5l=qO�˓��9��OL��p�¤@����ÎU�@���'s���ż���r`�^u�ȵBy̓q�Ex�g��H�6�&�q�I�z/�1�`bB
�az����:���g���~4 � ���b��܅�	�o�Q@�A�C��p��V7�uFy=�g}���k�&p��7t#�0�B��y�Ħ`��X"Ŋ��;+��������5�O�왆�4����S�P��\kW�'D
�&�� ֙�RN��>����Y�kk�lp�"O��:2�t��b-�i�}x��N����ߨzP
]�!K�.�f�AS���r�!��\�h�B.P?=���f/R�$���<��>��̛&�ZEd��#W!���h�<Y�'C�bx�#N2g�I�E�g}2�'�|�4���C�*�*�>%�8	+�@%~�O�q�7��TH�A��3,�8� @��y�LN��X[�옃^#|�
�H*K���)ғ�hO�S3*����c/�@�h�ĐB�	 8�v��EÐm�RxX��B�U&v��b�����9���;P�I�3a�#+���d"O6�h�@���%HFe[*�*��5�Z�OS�m{$��S�N�
�k��NVx�<y���N2а�SJ޾z������p�<aD��+F`���
�D��l���_a8��'�|�6��$%x��Z�~���m9}2�ij�{R!�4O��"^��r�S��p?a�O�<��� �8=iDKT�V�9�Q�;4�h����>4�L��(wu���3@l�'��Z�s����	�=ؠ$kd"����)1a4D�䪀EQ\4�diɺw1�\Y6.��L��	U�U;��O�X�<b�!�B�	''jkEg�E���lJ	sΞ ��l�z����g��*6��`��Dy��|Z5d��	M ��	Z!�Tx���N�<�h��7z����՜�ԥ�P��H�'Q�$:ʧ{Fh����#lqڅi����|Y�'Q�}2ț�~��쌼|,�h��Ǣ�0?�)O\��98�@� ���l�Xd� �'��'�ֹ�጖{1t���HF.�"�3�	d���)�BoY���]�Զt9�j�r�!���(&v2=�h�]�D�p�hZ6R�!�$� ��)饀��J��H�5G���Ox�h�&�Xt΀�v\�hjTI�sr�C#"O qq�i	(`�5�i�*b���G	�<qM>E��'�¤�RG��g�h!I��(�F�a�'�i`R�O-;��YC"�5S�|�Y�',qOƣ=��h����jO�y$:!ÓA�@�.݅�J�	�3��
D��Q����!��1�B�I&�B���
�)�z!ñ��Q�b��F{��4�+=��ŨĬģ%<"<�ř�y��I-�n�hQr y�U���hO���d��ZR@\he�̼"��'O�*~;!�ą��6���@Gc���[���"`$!��-�]Tn��v͞}"��1G!�0\���7g�pd�R�IڈVb!��p��dX�]m��1��<]TQ��E���%4%�eq��'[�"M��K��yR�Z:ox���^���d
c��y�♋~�R])�lQ[0X�N���=�Q� Q��R�*�j指�4eqe�Ƹo�6O��=�~
�CZ�n��F�yόH�d�G�]�DDxJ|b��GeOJ-h�&I�+ �{ �C�p8�L�q�ߞ{RD3a�!rQ��[��=ғ�hO����d���.1	������K�lB�	��!O��,O~���I]!j�ZB�	;�ɺ���T>�Y�B���B��ܟT�c9p6�z�U�',��g!D�4IaE+o�HQ�4�^! ?��{�- D�T���$N�|*saۑ5+�U(�K?D� �&��:�PDx�F���=�(*D���.֋
D�4gK�޾q1�n*D�x�1)�#?h5��ʷ<A��ʱL4D�� ���c�&6�"���*׀���"O\M+C�Բv�p	�#K�H'ZP��	QX�ĸ�ER�?ᶴk�eY�H;��"C;lOv� ��fC���EB��[�;�J5"cJ�>IH�̆�6�N�"�l�Wm�i��.�(F�����2}GKE���r� �C�E��ybb©>�h���X�c5���yH�#��A�T�
'?�]������y�#�xP��� h!���,ɸ�y�hğcY:U��B�2�x���G��'6ў�Omt��6�� >����V�8�Fx��'�dLѵkK�yXp�qn��B{��B���3O��@c�#v^����bx�p!4D�0�a�.ws~p�6ņ=ɬpB���O�u��ox�<S��8W���b�ƆV4~�L6D��JD�����(�49D,�5�0D�lq��Oa�=+���xN���0��@����	/� i�܊H�L�T���W�B�I:aN�A�u&M�C��z`�_�!dC�	�D�����EO=�vlv%�6y:�B�ɴkٸ�[�MX/�,��ԇ��
=:B��-�=�a���@� X���Y��C�Iai*쓦�*�Z8��;t޼C�(�Q,�y��-�P�hB�	<,.��ɥ.�5�����ϯ^�C��24�dP�O�x��X����B䉇;�d�0䔾!� �#
N �B�ɱ|��5�F+	���I�� �B�I:V��hf�L�<`H1ƅO�f3nB�	�-�N��6N�M�&$�2+�z�@B�I>KT˕A�5q�$�ʃ&V�i��C��$��,�"+�I�>!��� r��C�I�^����r��4���dB@�v��B�I�W���sv�32�0j�]�_d�B�ɸKd�BE�Tf�(mif�Ƴ�~B�28��9s��pd1�JE,�hB�	.)��+�V�TLFuZ���(�:B�ɩ\d�Y�#G?Z�vk� '`*XC䉝�d!��|�l]��Ԓ?tB�� =w��9W�+n�8e���"d�B�I5\�-�P&�&C�`���y\B�ɮB�pA����t"�p
�UmENB�I�{�,-X��ЖB2��q(�5i�0B�@M�<��兂I߰�k��QB�lB�	�~�PsnU$v5��6�͌	U�B䉙C ^ѫ�G�o����w��4&�C�I�H��M@҉��_��qv��.�C�I'����k�EbR�Ibt4�B�Ʌ3��P��T�+�� �
���B�882��&��t,����Λk �B�I�hH��� v��HI1�Z�AB�B�I�s(ٳ���3~�İ���.B�I�L�	���	�z�@��A^�,�B�I�+�yB�N\�
�JK��.�B䉝�0�`lJ,H.8��5��G�C䉷�l	h2�.#����
��b\pC�hҠ�����.�A�a�
6&,B�	�
�R�� iBSM�K5����B䉥G�P�*`�D4:��dn\,e�B�I�n����f��鉕IZ�C�B�I�7����D�g�މ(#�M�e{�C䉑T�:D*�d ,D��#K�6��C�ɚU3b�*�X֭���D�fC�I�(�x���o�����c��R�;��oVX�t�`
�1�0��� t$
���,R�H�X� ��E&�y�P"O�	�V�T�(�(-��m����E"O��k��V�.H9��m�"NZ�h�"O�HB�,
3/t��A8+(���P"O�E���B �����R"��p"O[!��?D:����λ-@���"OҤCu�]�s�*�S0W�h�|P�S"O�t���,b�-�G	�y�����"O&�1#�[g>���jG;����0"Ob����͆Z�:�{IZ0x�n1�u"OR	�壃�,1,	1 (�k���"O���`i�J�u"]�g��丒"O�袰��&{���
a�̂
*&(A"OL�ˇ]d�v��VÁ&( EX�"O�M���ϣ��yg��>uZ��"O���6 �E��`B��<�pը%"O�i�t��AS�(�'Z5�8<ф"O���G�&�Ȇ��#uh$�"O�
���`�*�ITC!wx�Ѫ�"O~ux%��#uJ�Ƣ�<k��P"O�9:���Yd�<x�BK�TY��"O2��F���zU��
f��*c��"O� !F��r��p�A�̧i��5�D"O�-0�O TP�yC��:F~�C"O��`g��2�H��")�1B�ɡ�"O�ȩ`��<#W� *FI]�,FR���"O �9�%�6�
�!m��j!�H:�"OR�h�-��Y-���\><|ٔ"O��J�EiX�f�ՓA`�J�"O
)Ro��E���%��t�S"O� ��6s����S'�y��Y�"O4V� �h4�	+�Hӓ_���"O&<RJ����Y2 ��5d����`"O��SB
5_��r0
�!��h��"O�����c��p��?H�Zq!�"O๒r��CLV=*Ɨ�v�\�"Oj�HfN��X�tc��%I�85+�"Ox�G��&_�X�8�D�Z���x�"O����_�a�&��B�K�
�ܔ20"Ob�H���=$	��ąE���"O��3P����TY��T1����"O� )e%�}�<�b�ˊ�Xd$ �F"O�9��-�Gr�@���:tW��8 "O��IsG��D�(�*AЕF1�i�g"OrP`&�C��X�[�F�:�N���"O�鋷e\���E�dK�,j�0t�e"O��[�	�(V0��A��!9��YbA"O"I�m�,�
�h�F��h9%"Oy@�C� `�@�j2��'s��"Ovp[�£S�2L�'��G���r"O,��Rf��k���r� [�Q�0!�"OXD�M�L�zp�6*C7x|h�"O  SgN�S��u����5� �"O��Aā��v�-�lƨ�
��G"O`Qyu��	/�t��
wMPmZ�"O�I�2��7'���
����qԘ|�J�� �a��OǄ}ؑ��K�.����F�]�'�(�ƭA;��������O�[
�d�N�D�N�7���ēR���Z �Q�l�d�L\T�HbR5�q�EP�2D�HZ ���'��2�V88%�Ä��>!
� z�@C���a���`2�B8���bL	B%�m;�IX}��2�|؀���5����`��y�m�2��p����J`Ti�V��ɡi�Ԙ��`@�˼eG�4�'j,	!q��LdA�4ȗ+�y
� �5K �h��x�!U���Qm_�Ǫ9�'w<
�Gv�g�ɸXr`� ���4�v�.k>�C��,>
|�D�J�P0X�͜*^�=�T�AI궐q!��5��ȡ�ŘJ�L��.K�<����Ov��A��G)n�`��R�͠&��x"ᓑ��a�g�5��ɜIњ8�5��
*$�]A�bM�G�B��Dɢ\����RB�5/�(`�J��H�Q�D���*<v=i��i���y��3}���.1������U�	��DWZr��I�:M�&�T{��f;���@����W���U_�p�#,�O��a�I�$n4��]F85�u%t�v�|��Tp"I�-,�����K�5a�.��#�����wt13�,�2}l��{�DK%�:��
�'�
��G��oA�|�Эh=��F�)x���
�3Z(l��	hhe �F����O"���@	s��9vg��<Q��9���1����VO�3GM�'h��S�AJ�O���h��s�Yچ�ѻW� �d���rh��P$n��k��*托o߈͋��#�"ק;#���H3 圀sS�V%8&��v��!Z�ѴIH�s�>h��┢`�0�倏�N��\h*Ç/*J-��I�J �T��Ɖ�c��0gk�%�v�O� �+ �b��T���ie��`V/�
w��1"��I&�q�F*}�����C0*�*��U���x���'.�2����q7��b�&£Iv6��B,p�C���.s`:���-:����?�SC!����ʌ)�C�+�;t ��+a�<��$�j���%*�/�.�����lCx�&�ٳ_�<���S,r������h���e�R.��'��%:k�PF�5PY~��	�5o�/�).�d��w�Q�nG����}u�E�K�<$x���$M#	KhH���P�Z(���c�'d��� ��W�� 0$ᚓC�����y�.q
�撘ps>��gT�#e�fP$fo&�I�烲Q}���ዀA:�D#ζd;�=�'�䝚w�!7��0��@&7 e�5�ߪ|�B*��LQ*S��Z����A�#4��4���<�λv�P��l�nDx���J�-��Ňȓf�޸�f�%�CU+����`3��͘4f�eYB޻T�����	��g�Аq�&�k�+���I;b���R��S���B���{����ę(r�l�#���<N��{��ʅ7,.�هf4$J��2�Z�l(S��yb"h� ��-��I��K��-��]б>��`� U;wLX��"H ��#@4�X����GZ�#7G�&%!="A�C�e�� T@U\00y�w�iZ����R��LU�U�Ӗ}��<����K&�<��F+V4�D*]�=4����$��d�BeA"I�������
	K,����.Z�4���|�����JR���A�'����'��%)���Ő�=|Ą�I�G���#g'p��OͶ��!8�D �
3D���	;��\�a�]E�ɐ���f x��sOM7���	�CY��K	+T� X�@dK�D�����j�d��(��p����Aʁu�N8z�"�[J��@���� p���R&�%��%�va�@��@�4@xѢ�O2`�c����p� -J7'l� ��đaB8�Շ�5*ے���d���@LSV���C��D�G-}ޜ	5E*}��O3_���}�'l=��.�J�" ����$%-O,!�  k����T�Yˬ�cd$�		q��|�J���lQv�ߔ9���UIH�K��q�Ng�a|2�´�4�Ȱ�]e��tr���.D�A�	��mIv̦4GT�I?���l�Nn���u3O���O]+�E9t˅<��۠�'8��tϚ'3jz�ڷ'@)�6��c��g=�Qr�&�m~B�ܪ�p`���|J|ڇK0Z��{��\���(��K]�'�t)�o�	w�0�'>���i�f�ĹqՈЫM�212@`
.�BHc�{"�t�s@�:m��1�G@?�(Ԫ�l�<��&��L� �6}��%�y�e�;1��!]��!�D�/(�L��
R ;'�-�mP�2�n�OJ�c��ڣo��i	�VI�{"k�6O��K �w���c�5��r�D2E�TRM�2[��Kr�J�}@��'!�L%;�%�>&R�$�L>E��J��3��I��Ӆ��N�J�?y oO	Y�(82h.�IR�.v ���1>F����iA�8��c~�\��SDs���$�J�x�p���+J/S�
A��IV�T���UL�)���P�(�>�b�!uin��S��e��Ju�&R
9��w�8("A�<��}��	�Q`,��=��DS(1ȸ�p$��f�!'�+}�'\���A���*�lT['*{�$��ȓgZ���[m�l��^!P��4�]���
��ڽ�ӧh���u+2*�Pd�@�|�mx�"Ob�"pN@���
���eA�(
A�>	E��ǚ�iD�4O|pKp�H�T088Př�>�~M{��'��am@�%Ϟe��E�h*��S�P�����l�f<���X��ys�M]��"�s�'̈�ZpjQ64[���|b��M�H���- �NC�m �	m�<y��l���qB�)Z��Ɔ�o}҈��]�r�|��I	%-\�՚6�7(cdX�/�-_�!�� f$k&΋�i�^
�։U��|;e�|�EV�T��x��ɤK�6�ː ��Kz<��,J�vbC�+��٪Ư^f4\���䇦THC�	%*�]c񂞏U|��0ǈ�K$�B�	�Nfp�ㅌÀɖ��T�
�1&�B䉔V�̈�J�5,�2M��f
��C��JL�Q�V\�18t5�@��0B��4M�^�"U�٥z��C��¡e�B��K���a��oZ��C�K�~F��!��D�?"�>�7�����,9iLA5#�C�(���r|&�Qs.ԟ�eP��J�BŔ�r~.�y#�T�0?�W�D��E4�Ī.1���bX]X�ܛ@��VZnd'^���w�<H
��r2GӽӒ�q�)D���⁤�&�bD� D��pG2�	
�7!�%���2rB�����"lC�DsV"O��S��Ê>y�ƀZ�F?�0�bhɻ�:�'�th1�E1�3��Y�)F�����ȠN����d\:v!�$�T�V�y��Pa&��D�7q��y���aGN��L?�����l����J�c�d�剘'��*�Nn-�����tDעe�R�z3 Ğp�bC�$�f���F\���)b$'�p��O$!cD�"K�������.\5��;��Tcl��;5!�ZVǾ�2p��>\��r��6��IU�+}� Y#m:bb?O���1낽TD���T+Q��EOdA���2�Ҡ�2!T?q/�8+�ǎ8}j=S�	-�O�$�qx��9�oߺj*��ȴ�'M��/u��9x>|��3�~�&�`Aͮj[!�łS�h&	����ԁ"c!��R3+>|`�F�|���y3��+SQ!�DN0�򰧊%]���e-K=!��%pr��r�jĀ>��4CD�E5<y!�K-Y���+�D�x�^�b�
�?
w!�X/*��tsD�cϠٱ�Ă$b!�݃aFPT�r�F�H���D"q���'����A�,z�jq$ ��>̔T�'р�@�Uo�l�+4�׊ �ҜC�'�R��6� �q{a���0�nYz�'�HD���N
`>)p�O> ��b�'e�5J,���I�%��~�B�
�'k�5�ffW4p>����m�z:�c�'��������~9Ć�&-��49�'%(��'�Zg�dB�ư����'��r�ڎA ��W�L�	R05�'�r�2�vݬI26���A�'�E�bB�4}��E�F��#	�'"���4F�,��	��'�,�� �'
�I#�hK�r�>X����k�Ɯ�	�'����a#���y�
�fȐA�'kŪ2�Ø�1"��4C�
8��'D�	p	ۑ	���(ڷ~<��	�'�D��5�D�T�XtX�d7i"�	�'}]�GǦ2�|x�NI.{c�b�'���3b��O��p!�*ڳ>T��'�.IZI�)�L��,"�@�S�'�H�����* ��lbv�O�&�xLK�'��q`㎎_ 	�N� �����'Y���u[ZF�ѧR�"�)��'9�����V|�I�+�zѐ�'�Z�H$ʜ;w��X�����>���'�D�� Fӵ��&�-<�$�4�3D�t��%�.ZL�!qg�F�0�0D�h��K%D�̴�Tk�yK�h�/D���
�nI8���K[���J`�*D�0B2MW�#��qS��E5c���r-'D�� ���a��D�|s�F=?�LBR"OH�pti��Yk��q*Ȯ?�HX�"O�=ҥD�9,VH���Q�.�$�I�"OLl#���)� �q����Y��(#�"O#hŷ` iP���g�12"O���q�ʗB�d����X�b��d"Op0A��'(���R���nȱk�"ON���l�%NLp)��$�#"OK�)��RP��.E�8�3����y�`ޒ:;ݣe��9a��GC'�y��-_�|��=e6h97���y��^�K�Ԫ�F�\�b��#  ��y2k�5�#��f�����y�C�-L-
9�� ��S�<\�B���yB#˻|����	���*���2�yңΕ(k y����d��Љ�I�y��)
H����Fh�PX�G�8�y�%�\�zI�S���h�pՁ�H���y�l��*�\ˠ�Y\�e:�@��yreB�d)84� �V��`pj����y"�DAH��2�
Ȍs:@����yr�
n��P��Opk����$�y���<邹ʗ�[�wu Y�
���yb�]�ľ�����<��Ͳ/���y3mB�Bf�7�.�-?.2X�ȓc�dX��ȂV8	�DX(<�
<�� E��S��JU9T� �.G&"����+�v銐$�V����O�
T�0���G:�2p�%$ظ��n��3���ȓNN��h6��a��0s2�$�N͆�uK<�{��	�5ߊ�����3�ȓmLR\0�-ɺ/��q���[�a}D�ȓcMlU�G���%�c�ջ"���D���9�׽f��$��4�$���uX"$@�̥x�<���lͲ_Lr)�ȓ<Q�3E'@:f��Z�&D�`��I�ȓC�RZ�Ɯ�Hނ���\$8� ؄ȓOӄ *1� -Q�d��L��.����r��xBH�&��Zܠz�����'�$��b �O�XA$$̔z�T�A�'|$b�@0�~�/Tr}�p�F%�y���~��-�Fa�8��=����y�K��Y�*a��g&3����jރ�y�	_=d�Ԡ��"�,#�4Q���
�yR��D�J� ��nҨ�Ee	�yb떀N�<;!�ҋM��Mb����y�B�%���E8�n�x�(*�y��&�����׳::�4JӁ�yB&�'F��Q����0� 	�1oY��y,�H�"T˕i�1�~��Qi�yB�J�0�iSL(C.��7Ş �y���-l���J�D1Z�<|b7+ȏ�y��¼PP��F*�(�d��!��y�H^H���V�2C ��#ݡ�y2O�'
ő1GD�Ai�]:�KJ�yR&� x$(��ǂ�nZ�K�!��y���Y6n�*�h�,jQ���V��y�9�d%���
�X��kA���y�ӻ�2� "l�N�4�)�,K��y�;Q�Y��%�.�ҧ������
��0|Z�KN���Zd��'������K�<a��\@8i6����q,U�ve�M��CC+���ē��RB��-�D�0nY<1���c�PyKS!� \�\!�D���"��
67��um�Ұ>� ��0e�7|H�'�+<�=+T�'nlİ�%����|h�\�|���ɡWZȸS��L� x�"#%D��eFK��8	˚"����"}2�җ0I�9�㏚�8��?�ڷ/ET��]��3g�4�!�)7D������u�j�ۿp�4=�b�U�F�]J/O���T J�Ѹ�����);5�ꈉ�f�+��	ʂ�g)5=Z�b@ɋ�ꌳ`�G*�:sCU,����{\����,��d�c�N�	^�ށj�\0y�����;; h�+��D!v[���'����B�~$2=��L�;~b��p/��\+�i�b�C8���%�ݎ|�1"U�.���b�2}rJ�{ZA���4��͐Q&\��I�T�(�%g�)��H?M�AR'.�u�C�	�y��=�#�PMyD��F�?n���7��c}�3
�M�T���Oc�ȷM�������hT��EPd��3 �Yh<��G��q~D�@��/2|��'�As� ig�T���D>U��d\P(�<~�8���I�&׆0���T����b�-4��Gt�L�b߅ԭ쀇��4�N��2��74"�y �d���K�9�ޔ���T�D>�c����O�*;���U�C�"ٳP&<O����	B�$� Of���1��I*`��	��k�x2E��O��d���z�,m��f�gx�<)���(�����jW.Hx�4�!*#�$W/Kp���ja�D�^��4	@�$²�
��D,b�]&�p/V� ���qK!�$ʅA�ɃgcH�Z ������*�@ $��=y7�I�%x�@�!�'D���82�O69�3�c�Iʆ$��27�qxc*� vw��+1E?D��qӉV��yr�����Y�5�z�h
�% gε9 M��XȔ�a�)�����uW�x�_�!�AR��W�!�09��B���0=yƋRg��kḫh��y8��0p*�x��gÑ�B8##K*a;v #�"5lw",!�oE�0�ay�M'd?�h���	�+b�qb�����'`�i"逓"��|J��9��ؐf��e�8	R�̥g�X�A2��'b^�Yc�ˌ�U�r��q�5$� ��� �f��P�?�89��B -�>��.F�-�I�sO�y+4�2�"�j��@ҟ�{�0�:���
�p��Qq���.-��K�"OX��`݄m��`�p��":F��R��J �m�֋��	�L$�q��*�L�t��k��t�@N�#4Z��'���ɚfs�1J�FU���i�ӓ8��c��
c���@����2\V,� 'F e�ܣn�@�C��>���j �N���x�I�
D�#�O
�ѓӭ\�O��/&Z��*�z̓^��z�B�8����&��$B�u�ХK�t,��M�N䈢B1$Ӓ��Sg�n����+�$�O�4#鞈�����h�>lT�=����)�����OC6@BȐA\����,m�*\s��Ō?��	���n��8�tU�W$F'~��ճ�H�u]֠�#I֗|Orl·�'R�\q�"N�"�~����l�ޔ"q�C ��1�HFhS0�k̫R�TQĂ� �x��6e��l�Ȩ
�'�f�bu��&�9�ՆC�idԈ+	ۓG��x8�l�N��E
�*>����$�gIL#3�O�}���c/O=YH� !�36��\�׫��;���'n����OV�|���?{~r��TA^*_aj1Pg`~�'���UcR|��ܬ�_�M��m�E��v��B�$A����%Yږ��7�1}�ھN���}�'�^�*#�	AVrdp�o��sa�)O I��T���Hĭ�'��ՠ7␔q���y�+�-Z�j9		��:�$�0A���E��/u�����O��M2`*[�>��x��W�W� �m\$����c�M'0mp�A�� @���Md��j�J��yrF\̉�h_+	x.���?��?�0�\	.��� l���z`f�%�T��Gb�:��nIؽ"�D ��S⓭kl)I�٤~��I��]��?A�ĉb��-�w#�I�:<�F���9���j�Fْy� ��C(�a��h��d� �
4ض���6�na�'F�5c��I�μ�E�^�c��S�O�Be�p�ݵ_C��Y���>6+8�
�'�&M;���YMlY(��$��!-2}r���6D�!�g�O�T ��mܓS:� $K���<�/H�"��[	��>�,p�(QR$Vк1b�4$��q��B���"E�'XkB�Xw�)�'V.���R!�9m?�0Љ��Z���D���S��(t� g�9��iR��'{Dj�{B윐0X�'���(�d8"d�<��	��2��րӛ\�p,��M�\���7��p�c��S�IW,0hV0�j�n�Xp�	�`��2e 6�����'I Xx��ܒ\�̉��&$�Jѣ�{%��g��UI"��d�;R�S�`��?Ya$+���1 媌'^3PLi��?D�dC�-�%<Tl;�b3)��}js쫟�k٢��U�՟>E��(ٻe��L� AM�i)���F�̅�yªGz�|8�H_ڤ���d`7}�A.h�^Y+B�[S�8���?���c�CQP��s�:�O�L�f�Z�WL��׊G��yf-
�T�t}
���x
� Ƭ�G�[�\��8g���q��1�5��*���Ł[�r�1�:�X��ڐO�4�Q �L��hs"O���b �	\�`,ddٔX��X��ה�$�"}*�l���XL�A��<`ĭ[QL�w�<q��j]3p'V8+6Vp#c�^i�	8*4Rx3s�'�P���b �����,S��<H�'Q\��7��[3�=c��ċ<W�y��'",� �O����2�DZ�N�hI�'�\]��ʬqL���M��C-0I	�'I� y2(	?)���Ud�+O�x��'5~��@���2��[�M�*��u�
�'�p*B�!�1&h��s�'J�"��e��	X��$�����d�Q�M��G��OH!ӵ��^OF䳱��a48	�wO�4���ڨ�8l0#�ޟ=� 1�уy��z�#�O�)R��r�|�P�P0!~R��'��%�AP�c/F��'"�e�fg͍.���r1�M�GR�@��']�c��X}|�P�� :9D�J<1��qx(,�t�+�'knX�0���9�2�(�#	�*���ȓ<�vI�G�ϊs�v���Z�k�ܨC����5f�.!؉�L<I�"�(t{6$ӄg��h��OH<�����b�'�r�dQ*"n@�;$��A阢5x�����2�XpIŨ��xT� �ay�*�= ����EyB�H��jgfU�X�R�y�Z�y�e��f�!�^�($8}@���-�ē?UDP� �T��u��)�C�)���1\%Ne2g��K!�D�A��YJc�O����4IL�r�J�0�8}�)ҙ!�\c?OP�b��� -6�H��N�R��UO|�IdL��f���!�ZX����F��}K�
.�O�Ác�n�{��A��^�Rv�'��5K�`O��O=HQ�x M�"�@�HFMQ9e!�D4z������e��0W���3!�ܫ�v����Y�_P��ϕ*�!���؎���mY�Nf�P"
M�i�!�##r(� �+��q ��!�!�d�
*��b(��+4��_�!�dE�E�0�S��*�*� U�5,�!��%R��J��M����.ؿE�!�$��
����D��ܛ���\ !�� k@Ѐ�c���p�t��5!��7�r�j���2�$��6y!򤌳c&@=��+E;��T�%��7!��\h� ��Ȕ�v=|�R��4<#!��DF�h,q$�H"z1��)_I!�X�ID�ȃN	Hف���-xO!�dƈc��#� F�5���$�C6g!����yY���T+�R@��"Of	��J@mj�l�Yy�"OP��rCվfju���ẅ�p"O�E
	
Y(�� ״e߸}�q"O(X$���	d�so٥?� ���"Ot���MA�y0Y��Y�f�Nh@�"O��"ݠ	3����۩5�<��C"O����L�Z�T3�k\� da"OȘQ0��,"6���:]�(t��"O��DF·a���P�Eߙqv�#"O���r�[�m�AS C�gM�Qe"OxrD:@81Dר �����"O�%�C�[ x���& ���"ON ɕlP�TP(rgÇ&+�>�Jb"O���-�Ir89���>/	��@t"O��� m�QYF@�̣j��� �"O\��EɎE�\�dd޺B���7"O2Ő�C�afI�0l�23<�1�"O� V,R���QL`t��ޖd#
QY�"O6�� EL�|0"��I�0�� �"O�EI[�Q�@i��N3f��%P�"O�Y��@1*�dɘ��'RN�$��"O0�p�gK�m�ʩ:1.��r7p�"O�%s5�Y2F��Ze�L����B"O��{��Q fहG��]�z���"O&TQU��(h�p�&�j����R����6`��iRX������ a�Aqi�c�tʝ&v\$,�9�.�P�]3�M�Ԯ�%R\;�"����s�f�6*U�h�4BF�ga��pA�h�Pрƀ���)��c��/�=��a�3L,�q` ̱0�^H�”��~r�σ�0|Ů	�u	RY����N)~�Gk��Q��'�P�Z����0|���^�
�ވ��!
�'���Bw~"��tN���eIE���L�<�у*���ur��`��6m�'={RA�� � N/tէȟ x���ǉc	N���Eٛ5�=�r�79�z�0���?I]�恆=�?E�d�J���bf0��s�
��b\d��䕎f��+1h��7��l!���(H\��Oo�2|�##+!rE�!��95�ȥ9��>3e�$S��[��8a���">R�(��ޒV ɨ�&�4`.�%��B��ƪA���@�\>�S�ľi:F��+�&T�\H!�܏Z0�+M<�RI8�b8�G�O��\���Z�2��(�!~X�¬OZ�B��ԭ@!�O�>a�5�߽�t�	�&��+�u�s#e�$��� ڮ5�ВO�?m��꓆0��Y�%W����*2"�8�<m3.�u^���)�'Wd4)EM�k�Ѣ��)�J�m�A�R1(���'V����fȘ�NRm�Oʜ��O�"|�S��~Z���6"ހ% $��c�V�	�.IH}A�	���=��	SI��#-�?*���;�j�2�Ҡ!B�bӦ��W�5u�\�O�?�#ú4�+�'1E�,���\�132�cQC0B��	.��|�� ��M�C5���"�H"?��@׬����Dh5z��9�b⓽{�֐ a��aW ɂQ*PS 7� �T�� <�iݭ���h8wlT1����b䍩&K����� Y�创SLqO哒? ,���S�`��2�4�дi�",#���(B�L+1�сM��,�"�^,S�>�|Q���wk�,X�� 8�]74��劏x��͊M>E��',���M�B�C�n� /Cv� �']|a�1@P*ɨ�"֜-|:x�'�t��i	*N��Y��)���V���'#�	�DW���	[�3*'L��'�,�hq���P�D�!�JA=%�xP��'��0�J�5���2Wf�x�p
�'�rP;�Aŭ�ꅊ�)tf��'���2��t[���b�l�$(��'�|�YGb�2wZ��9�OH�ij�5j�'�HM�q,_M��ɡ�`͛d����'S����D�RCtU9'$�X�ܥ�
�'� Dp�{D�bV�B3Tt%
�'e��1���Q�E�!M0z��
�'	�	���_mA�q�`NZ�\iԈ�	�'�t���O� $��cP��*_ 2�y	�'�z�Hu����@B �Q"H5)	�'hh(��*�0hUb�"�؈��'�:087凚p����]���'������W�M�f�s�a�8W��T��'m�f$��d��s�� U>�)�'G�˖)欕�q"�%U����'�%�S���s椰9���)ZD��
�'��0�%��c�>e������E*
�'��-A��b�"��� Q!E� �	�'�^}S$����Q �k,G��L8�'[����l%�����O`xa��'���7B�$$?}1�i��Nf��
�'�(�"K	�pl1MB����
�'�ntx�.�#9��Y�*��7F���'q�8 �eA�#ޔ�
��D����'E�-�c����H�����r�B���'V�!�R�8oB��H_��r��>D�� �p�E�X�$\0��¿Jˌ4��"O��#�b��pXO�S� (a�"O��!Ƈq�4���;'t���"Od٦g��B����Ǖa��q�"OpQC�ۆ:D��U!ި]_"��"OZ�SV�սd򞀹�/W�-��)h"O� ��'Ƶ���V�|�[�"O�5�ʉh�VQ�6�(�0�"O�l�֡ȵK�u����R��rg"O���'�p�R��� �4��}	"O�P�Vh�:L�4E#0Ȼf�p8�"O���Ɇ>�|؊LU+_�Dux�"O�p��֊;\v�Y�Ȁ�*��5�"O!Cb�I�--���#�A��K�"Oh��q�c�<yȇ��T����"O��b
��~�4���ݕ ����4"O���ɾ�
s���%�U"Of<
��J� ��Qj1��(9d"Ov%����n�z�M���%����yi�2���@$�^�r�[���y©�i�u�e��U5<�{f��ybJֳJ�|�0�ώL�~,�P��y��Ä����/�Q�<`5��8�yb��/ 	����Ȓ^N.	:F��y��\�&<9��'\���t�Q��y�  �f �-��팚X�(a1�\��y�"��2��=��0O�T�Ҋ<�yMK���9��qn�P���yRe�#}�v)b��W�>�1"����y�]�{g0��.�C��j���y�ܭR�����W0B3��J҈T��yR�C&�����8^pբq�@��y��>R`���!�0}Z��͖��y�G E����)!1(� �"����y"�F���@ @�X-���[!�y�O� l���@�E: �$�yB�U�[=Z�b��Ǻ�����P��yҁK�C ������ȓe���y2J��C.):Պ׬=�(�'N��y���4�:�k��G*e{���<�ybkb��1�'�V1��Ͳ�y�F9�&�CA͚ejfj4.�y�!�:�c��� dm6	P4���y�`W(�|�Q�lT�Gr�� �3�ybm�3g�l+1�څGp��A���y���i�@�C	�9fDP��O��y"h���@�[�#�>�}S�j�y�"��{�x`�M;K^쌛�
�yr���\�� �īG:U��`�;�y�7z�^�IR�G	�-:����y�B}�d�x��B(D"��$��y�ļt�jihA���o��a�A���y��-�ycd�R����Q�х�y�W�Dm(��� Ui�a	��yJ�x̩��� �vreI�KM��y"mX9�e�a�fo ]sA��>�y��O�B.*�{v�[�do&y*T�س�yB���t��D�/`L�(d���y¢\�Z9��0R��@ܴ��T�G��y��ó�ld����I�<r�ь�yb��g�L���N�&�3�aY��y��^�q��K�(A���ү��yOH 9�8P����:c�0����yB��7?hJ�Ц'�"6g��JU����y
� JQ0�a�:m~0 ���%|��4�"OZ��U�{�8`Ad&�`���c"O�x×�V\W  т�;t�0��"O$��$.�P���膕6���[e"O䌊UB�GQ`�k7I��U��9�"O�h�&�pCP�1N� w;6�Ѕ"O��Xh�"VL��9��";$�p0�"O�ݙp� p�`� m�S<0Ÿ�"Odh��g�3.�H���p�h�c"OB��l�	(|Zab�%��|�:��a"O,$���įO�p�(t*݆�:Q(�"O �5���(P: K�(U׼�'"O�<������ԑ�L�K�~T��"O�yr���YX~q���T��2u"OX=��[�]R�HZ�D��<ҧ"O���V��\����u�V.u7"E��"O��k� H7������ȗh6���4"O�P���	Ăݓ��#D��e"Or�����Jd"��������t�"O��C�Q-עa�w܏q�`��"O��%��(�V%�����\��L%D����͝-P��rI֮�X�#D������'H%bTa�È7װpra�!D�\���! �e��+l��v>D�pADH .r�b�G�{Dr��e�(D��(��/#�3s���+К��Q�1D��h�&�|�C5ȏ1g�,@,D�\Y��ӟ���Z����%h� B@�(D� �b���d���H '���0��&D���Dπ�
G���2%ې9k����'2D�@�GQ�-��0ʄ�[``��3D�4Xa�[�c����J� �3g7D�`8��b�4`a`)� `M��rA:D����9+z�)s��5⚵부3D�t��߾\�Ph$-��n�r¥3D��镈G�2��|������I�K-D����ޑ�L:enR��~t��,D�4ه^5Π`�v9�U>D��C-�2	�ThP �S�Z��/D���U��lL���^Fv��u�7D�q��9m�d�Rӡ�qK�y��*D�D@Ԏ��hu�M��@��'D���gII�,#�A�1OF17,�cb�$D�7��^��L��ϑ6���"�F D�l�v"U2�=����)/���Ei>D��RbZ�GQn���a�8M��!D�T�Pe��5
de�w��nB&t
1f%D���ޭFN���#K��Y?��E(D����,��`xL7f9���w�$D�$jӪ�����%��R���n.D�(�E�Tk��)v�ɺ1TA�wf+D�t����hD�-Ҁ�ǵ�V�*ï5D� ��g�
TBԐ��qB���5D��B�;>v!��F�j�q۠$/D���e Z8��X�`iIim�f!D�xs��Ιm���f@4V����-*D�0&ű!�j�:@��7�̠@PM'D�@��"��4�2vC�q��D3D�D���3����J��$jǦ=D����^�&<Z���#�k"�;D�� W.��{
�M����fD�sU�9D���@Jض9����̀�0x�l��7D�p�5�*0����`������%+2D��Qg�˂o:T}!�&0e�`e�#D�� p Sw�Թ@��x�슙_X����"O��X`%A+j�)��N�]H"-2c"O�4S Muز��0���&��"O
��ġZ��[P/�c%�iy�"O��I�$�m��z�`�yB��F"Oj�z%��p�@��w��1"O�<�#j�
f��i�%Ͷ	j�"O�%�ːE! T�pj�,#�֥ �"O�,�L�\�N�i�"B�V-�B"O��P�-��cPB�q	�l�*Q0�"O��R����e<�FP���	�"O*l@��Jr��T�ϙf����"On�i��͚z���#�ĚP�`�+f"O��{���;u)jhy�+¾���b"O�E[�Y=x���)�$�X	��"O����"�"jS*tIA�	Av��V"O`���^�#��� �'�?pղ4"O|��A+��Y�ҩ@��ϛti��"O�M봬	1����QA�US4"O�{�HL�l��0��_�(��"O�|B��;?��ꃦǿBQ@�{�"O�����Dr<���VMXqi�"OvL:��4
l��S��](�  "OH�r��B�+֍5oY�>�i�"O��h��X;}1J��q��J"8F"O�0ن�X#~@
0 �jL#+C
��"Old[�9a�4ab0��)6x��s"O��A��9V5��;����-$V�S�"O2��vC�b�~	�"�4`��"O
�7Y1j�ѐ+
�x�|3b"O<�`T�K�v8j���8F\l�v"O�As$�	�P�07�v߀Q"O4���S�O�9�R�S�&#���g"O�)(1I��3	���D��'R�:"O�7j�w|LM���(1BŒ&"O<ႈ��{���	D`�dzpu�B"O.�� � �&�����VAh��"O�Q�   ��   z
  �  d  �%  O.  #8  �C  �O  d[  g  �r  �~  &�  ��  ��  U�  {�  w�  ��  ��  ��  ��  !�  g�  ��  ��  >�  }�  �  � � | �$ C+ �1 �7 ,> mD �J �P tW �] Gd k �q �x �� <� 7� -� �� � .� �� F� �  `� u�	����ZviC�'ln\�0�Iz+����K*(ac�
�bڴJ���|��ƟH�U�>�D9 L�BpI(��
0���3���%m�������D����p���u'���%��֖9���o3 �����Vp��)�掔�C��dʃ(�.g�^�r��Y�: �rÁ�c	 �]
bo���S��`Pe��w��H��%?G�8Cq��S��U#�M��?ɇ�P�B��L�Re��Q���5���'wb�'#�+3_� `!�iN	My�p8C ;���'�bo�rʓ�?q��Ŧ�����?iԍ� X��&X�F,lp�!��?���#c�'2DL�G�'�>��޴�~��O��Q�S-Ѝ:�ư�1!�7J�� ��'��d>8L�D�bY�YS� �!�2˓�S�N<j��F����i�a�;=�괒5��+f,�睯]7��;2�J�2a�%N�z����O����O*���O��$�O ��#�S�G�g����ѷf��c'�ȟD0�4U��d���'6�7M�ߦq;ٴuC�&�' �D{ca�*3(i{7-��B��P��,�7f�?�Q�ke�6��r`�*Lm��� a��mח+�0�R��O�Lm��M��'��T����j�Z ˕e(���u��<\\ѫ��;��&�US�ic��z�b!.�\iy�憏S@�Dk�oh�
�n���M3�/�:�>��,k���p���<,���� ����i��7�>d�j�Q H�D�l�;RÑ/5��\a֯ۄ2{=��߱ w���D"[�,�eb��M1X�:5Ap�^��rڴ���N�o%�P��-R�q�a`Q�ğ=~�ģ�A�x��t��C(Ԡ�w�^<�2H�	x�����c�#5��@�	�O����e���*��x�G]�> �e��Zݟ�?���?�e��"|���'Zr!��]+^@�5O�On�����D$s ��'�"8�$�'�6���)6��_0|�FHI?c-P�Ҷ�Zw�&��Ȝ�c<P�s"� -e�ax%؄D�p�����Kk���G���m�R�LU,���g�)��@��'a����?Q�OP��@�u�N�;�R���I�'�"�'��OQ>:��>�F*�P7��q�$0�O����H��	*��Ik
��H�
�bS��<�I!Jo�"|қwj
ɠ�B�;v0��s���'�B�QbkG}��:��+mh\
�'z�����|6iנW`� �X
�'�X��� �q�X�A���h����	�'�J��`ʋyk���ʆ7!���'���Z��=K�$
���/ ���
�-Dx��i6>�2�{1��]���cFJ6++�C�I�+XL� BF�'a�d�6AE
]��B�	�d�rA�艌^��HJ�A�@�C�	m:�3U�p �քF�ӷl.D�����cEt�0dg?aI��{ł6D�8h�ǃ�Tu:$��W~TF�I	�<g��G8���pK�:n�8�P�ɦM��]yUj;D�(�.�q!�4�Pm;O����L;D���芢V��M+e�m.D�b1�#D���$��C�ڀY�d&}"�KT D��ۤ&�H������@�?<O�{=O�P���!X��qb�lI~������$8�FH��j�~�I%E��yB�7y$�}h��9�r��Q2'�TI3�	-���=F#�erP�ڸt��� ��/Tax����?���?���k��O؉|,,�B��]%;/�E(O���2�)ʧV5��iاU�����^OU����I �?Y�A �(~�JdL#��@2�C����?�A\�O��N��-c&�A�
��~x��)�fȼ�!��1	$�h�۶4���PD�m�!�$Y�2Rhy��!��Tyn����/�!�YyI���G�@o�fb:�	�4"O����/�X���quhZ7I�C�"O�����6��ቚP�xa�U&�MS��?��:��)[3�S��?y��?!��Ϳks#�P阹�%hT>k�y�A��'(v���',����j�=s&\[P)��&�j-C�yb�I	��y����H�d�$��@��@��?��O���'�1�b�'�2HC�U
�cT�C"���'��P�!�p��H�.�17ȍp@m W�HA��4�$��<!s�գ�.Q�h���ѕM�T)$�u�X��n¾T�&��<&�صoz#~h0��*�H��۩���A�Iфpp9s3� G�C�	���l�6��m(�L�PI�$_E��m�Oȝ��I&T����לKK.�c��$@B�I�=�JR�8�S�gMl���$�����%$�8X/����	�O����m�hg�$Y��Bp��ل��O�$�&~�4�$�O���Y,؃ď�`JZ@��� �M� �i� CV�O1��C���6gEx�(c�'�̴�k�bI�
�MJ�W�F6m޶M���g�V���P�ե�A�ax�(E��?9����D��%�*AI�]���*��B�F'�'���'�zq���^�|�p �R9h�P��pt�/:'�xqj'K�{r2L�tN���?�(O���ӎ�����	ܟėOm����'C�D*W=SrX{u-Ч}y�1"g�'��a�-d�D�b5"E?F�>�T>��O>r��#�X<1��c�&�,ZF	9�O��EM	7xR �K�fJ�}"S��:�xT���;aҢ[F~B+7�?i���'��O͈�;�����0�@����ک�H>����0=�����)S�IH�B�6��x2SD�G�'X�}����2uV�y�uE�;V~��sÞ?�Ms���?��0�8{�l���?!���?����y��ځ3�v2��|!�q�q�\��'b*��
ӓ5�6M �L�*l��S�@
5���<I6�R��T��*4�����_(c��ؙ���O��D�O�:fh�O�c>���dN�"��]jA�јs��p(�-�y�g������9gހ�`����D�w�����'��ɰHE�tY�ơj$e�@ �uJ\�+�lM�7�`,��؟�����dQ�����a>�E`Ů*]��2��]0��ꗁ��2�=����2:�Y�&��vx�p���=��թ""�Fɺ��H����¬��Fb@H�k�kx���¬�_>����^d���
<5�����O`���O���?A�r�D�O�Brň&s�d�Q��X�Lk!� �5Ъ%���7�� ��b�
X �'e7�O�ʓ5(	��X?���%��q '��di �a�� �=�<���؟�D	�؟��	�|�ҡܤw�`0P�MH��|��GԆP-P��2e�L�p��MT��x���> D�g(��yB�Á�����蠓�$* @3�S>btiW����O.�P1�'
�P��KSr��CG����˘WA�'-a|"fWsM$(ѐ��رɴ�ޭ��?���'m�\�e�S���I�
B�>�C����_$S
�$�O0��%�r�\���Br�(��y��N>�v��g�� ��4�LEʣn�Lv2aZ�ʧ��)ɳ6�^����J�F�#"E3���!�1KD�'vi^�p��)δ2��%����w��Q��E8��	�����O�}��'� �ba&��P�̠��̞&��K�<`��Ut:�팥[��U+�o�a�'��}��߯'�E1m�h`JH����M����?�q��p�2(M��?)��?���yG�6�\�pɛ�!�VD�BnԸ�y@�FƘ?�N7��Q4=&��B�~�Z0��B�?
!m�F��T���DF8�mZ��~�Z�*=�3�I���ݣ#�+D��DɡM���0?��C�쟴����h�?WDĆ$Ki!1�P�$$�KRb�8�yBa_2��P��=" ��z��>���R���T�'v�I�[�n����4%����"	ǄTP�l��x�	̟�I���[w���'%�	��#ߴ�.p��"M �8�<+�BO�Е�$$J��p=�a`	 mC�-
�h t���փ�P2.I�ǢҪd��dM"\O����ϖ�?�ճҪ�P��4�r�zӺ�l�b��"&�< ���e2ق�ߎ17
�A�"OV����M���9��Ytxȵ�|�A�>1,O�H�%��e�	�g(	�;@�Wy��s�ٟ���*Q�$,�I���'+w�5;VH�B�>q0��!�[-Fˢ��#��&p�LI��	�9���ˍ}��P(Lh��^"uR䐘a��<�0<IqB���X��ß��	)_[���s�ƶS�4aj�s���'����S�&s�0;�c7Z|�2ՁH������ҟX+# F<*o����XpFx��F�O�ʓ}4��iR�'D��p��8�	wh����}�h-�	� �֟|�	�\���0�GJ	b�x4�K��?�O��4<2�dx��ҍG�ʠ0#���D��:�&@a�Z�Ea��h��yP�i�%`�h�d�/�
5K$���hт�O����O2�d$§8�05;s����
uKE�<m ��'�\�	y�� !�.�]��!�BY�Qլq���*�ko�>I�� ?*���s��,B<EP�<O���O���^&2�P�����O����O��i�-��O�5:��딁ףD�8�z��C�Y�᪰���Nm��B$�N�@��b>}3O<��Z�(9T�6V�B� �"�2�VжG	qV&h�tLG�@�|◩ڗuG2��C����BQ���%�֚s��	a~�+X-�?A��hOlmS�o�)6��%H�]�n���&,D�@�!�G��4D�!@��v̖��w�<)��i>���ty�eZ�5�h !/?l���v�U)��Q����'���'9�)a�����$ϧV��v�īV��y�J�gD#D�
V� [��Ȁ�S5f.uӑ��'5� ��%�Vi®�C�ʉ(*�H�� څzѠU�tk�$D�V�!KL�?zD]���I)
�<"�&�kl�i2^'l�jȨE��O��*��O��;�g<=����۾$,��I�"O�E���t�%�T81�µh2�|�dkӎ���<9s�,&Z�	��g�D�,���Cp�(-�ᒦiL�D�I�v�~@�Iퟔϧ�nHC4�GD�lʆ�b�C�"�p3��?�>��	:->�H�}�(�3~+��h3�<B�x( �(R��0<Qፅן��	���	�
~�X��ύ���x��J�&��'Cr���]�ԭ#����0��Թ=������ǟ왠�ř����_/r���F�O��ft�����?Y������6C��7/�4��T�W�ʵ!⌞�Ln��'��)؆I� 2�$	��@@A}*���'X乡E������c��ipt-�'MX!�4B�R���S�.�'	�<�`I�1D0�����,�,�'d�`r��?���ih�L(aB�7u����Y�
L]:��+D���@��X� V\�q =�`��>��F̖=buR�j�^���b^ܦ��	�x�	32�"s2���|����p�����n	�@H�K�$k�,բ��v̓J��]��	���AX�~&|�Bd|�c�p�@L.LOz!+�4t�4�f�W$�>0�'5��' z�A��'�1����|J�� �Ŋuip������C�z�<��FE!]!.�!��K�R��CL\y2h;��|�����S8~����P��p�X��� jr�l��?O�����J�@�� �.]�p�3�!K�v>#�ĂV}L ��(ˢ7v|t���k�'g�˰jG
q,%�2�P \+�2�V�#�6�`�\�¡��D�7+����j��OX}0B��S���p0˟�ɴ���d�<2�Of�pS��@��j&͇�x�"O���0��Uq�$�]��ҽ⣛|�ab�ޓO�욖8O��1�B<Yg�ߴj���ElˁE�)��	��nUkq��4[?���TCULdH��Ɠ]�V[0��F�
�������OP��,�
8P��'�'�&��d�� r�D��l��[��Bv�ݵ���/آ�ት7BH�$*�I�d��[��%*��w%ׅ͊C�I�Wʔ`8�NZ[F��sT� {4������88_�qɄ�0��"$��/G�$�O��+U?O0�}��'i8a2aP�v)tHqj�;F�T��O�Tq��Ԩ^�&a�t�,�*D�U�'$�ΠB��*Tղ!�d��X����'�t�bW�δ
�0)�#�cM�Pl�}�t�ȟڍ0�H�X9���W�_�6q������(��/�O�b�"|*�c�2'��Ģ�+�2��5��	�q�<��J�%��E@�$ϏY���jl�'�h�}Z� ؽA���e5-;r��3���'�0�!ms��G|�������%�L�a�v�Ha4M.�Y)\�o��TPeIG�fj����*����d$���y8��(�J��∕!t(�=a��7g� ���)W�\ �>O�t���$m�n%�C�u	�#��Du�'���S��0+v�'F�p!3D�8[bnE,`��8�e��\�>�`̰<��i>�$�p*��S��=��h��6\*�C���	q������_�V)��cX�I��؋��0m�� ���[	r_���7D�X������	<r��
�!^�Xc8u��D�:Gy�R����+f�]>O Na���'B�r��	�Sn�|1��a���Ł���X1N�O�C�I�����7LH�x�LY�E#*B�ɫtOa���ޯ5m�����GJ+��O\)n�O��:W��IM~ M�$��2a��|���嗋�0<���(X��l�ӎ|8�&� ���u�V������F��n@l=pc�	>���%6�N�"�-̂R�V!���+p�~0b���#p� Zb�E�(�Z}7n*�l��]�	y̓Y���z���d�TS`H��;�H�ȓ2"��CbMƗi��3��C�d� ���	%�?���S�"tаu��,o>|����a�ɤc��Ic�O��D�t�r9�&"�:,�����	F����B4�d�ݗEM,��ȑ7'��)��DeӁ񒠢B⛦QF�E��
��d,{ǌ��c.�L�ss���mT����F08��S�o�y`S E5h�6����1��iԴ}��]�S�O�L��2Ś�}�]���ڲ%��e�<)Cͅ�$�`�8�����|�7��K�'�l�}Zc�.J�&hY�!
j��DYb���&�0�+n��F|b
�L��D�.FB�٨��@�:���TO ��bdi�����H���De1��ŃTV9��8�X�#�dŶ���&[7�� Hн]����i]&4.V�C<O� ���,\���2��[-�d���$�[)R�'��b���+r��pa_B4z�'�^(�䨉� 2(`��BV��0,O�5Gz�O-�'�{��	�j$�� ��H�Q�"TP"Eׅ�y��'��dXC��7_�调� �Hw�4��%TX5Jf� "Xn��!χu�#?�0,\+Z��@�"Uw�J��=,�(9ƫ�6@]���6A�6B܋�/�Z�h�Fx2Y��鹖fJ!,��tCef�h�jQ���x�)ߧ�$4p��6+��3�ʁ,�y��8r��bU+��GTQXĭƃ��8����|�aӧ�y��L��73˴�Ѕͼ�dX�:O6%8�#��%859�ϹC�h�`L�.ihd�F
%-G��bč��TG~RO],`@h�����4	�T(4���	db�
s�aj�n�0 Cd�0M�yU�-Q��Dʹ%���d͢Z�<Ze.T�Cj>5B�cW�!���L~١�&�@����#
���r��Oji��/,f����i� +F�k �|N�y��S�<y�®.`���^=!��T� ��F~
�HB�G�d�����b?E4#ӥ�\��'�[���<?IE�	�&Ƞ��T�q�ܓ�e��C����AB�H���D&Y)���W(9Z@���	����ą�Pv����;R.p�{�MW�v�`�%�
��<B���i�AN�TU�ȴJj��'$�X��>�rOH�$0X�Zc�[�~�lȘ��Ox9����P�OCd���$�6޼(��O�'@��DH�"OD���=H�����\�
�"O��R��8�1�G��ԂI!"OfQ����#�����2���"Of�zC�G?��	�t��*c���Jg"O H�"d{�.�!4H|��U�R�x@�i/�O��WI�?�Qx�fɺ���p`"O:�2$N�� ����tH$6ۋυ�yJ��U�F%�@|B��f�I�ybN �3�~����8C6q���_��y�"Ft�2�H
�|�0�,���>�6�~?QDKɅrP� u-
�|�� ���s�<�A,ɗC)�% Uk�uL��Dp�<�┾\3Av@e�`9��e�<�bj=g6:!@ň�>s�\QT,N]�<wD�	K@4�2L̑(�2Ks�<�P�g�X�2TD��JDhЎs�'3�iP�����k�K'Ɍ�F, ���`���!�)�I9zI:�0�M� l�!��?P��Y��EH�L��b��:�!��B69K4Uh7�ζfhʥa
�i�!���J�h�d� \U�ѓFH+/�!�L�Q���b���.=KrapĥU�?�B ��O?�r@)�ֵȒ��_LH�2a�q�<��ϵ'MơxS��=n�Q�k�<�Fl����ʖ�L���3��|�<�7ȏb&yJw���vB��^�<qb"�y~�I���P.��C u�!��m�l��)��HT��fmJ���	�����Ëi�.8�`��N�L��K0N9!��"7(�H3oէo�U����+!�[-z��
wa,-�t�ʕ$]�!��q�l�U�����{	�!򄜻u&�r1NC
e�-���_�}��}j�4�~R΀?G{e��h׶`2�kbڿ�yb@ӱ`���X lD�-�~�Z���y��[�=��=�(\�$%��
Eg�$�y��X>: ���O��!3}ѣ�í�y�@^Gg������(�ib�J	�y��
cjq�G�ϳ~e����� ��hO,���S&N��� C��� X�d'T1�C�	�ڭ�f��f���{��֬^�fC�ɎBp�aUiēe��(��)`NC�)� ��񒋀�9_�&�-+��R�"OJ��4x	)�4���R"O��[CK���,�'��=m����%�'K�������>�-��
��� �d'N�A��ȇ�R���u�ʖ������ߔ;nЅ�7A���� bd�p�z��5��0by�1�M�[0*`�`�J�6���N%;�'\%O�
E�@F1��]��k���UP:n��-2���.L��<�'Fg8�L�dH1@�83��
�r�B��%0D� vӚ~3V�P�DlhwN;D��r�	�4�l}���G,&v�H��,D��{��)�F$�(H�u�r庴�,D��Xc��"se��i�m�~��!G�%�Ol�ڰ�O�+/I<4�� ��d1X��"O�q��j,�8M��"Dp��y�&"Ov<���VH�F�� ��� �"O�ai��\�.Bl
Ŀ�o��u�"O
�3U���.R���Ɇ5S@��"O��j����1���B���|6$���#^$�~���]O�j�5-D�-�M� �W]�<�CgU�o����g�Y ,�q��`�<�ūΠs�.�"��/,���yǢ`�<���ގ$v��P`��N�Z�vW]�<y��X�okP�#��N�aT��[��Y�<��Ј=	��Q��^�g�ܤ�'Ξҟp#d�&�S�O#�љ�E&�+��D.*Ξ	��"O�LS�J�ֈ२�-^�x#"O�$سj��B��EV)h� a�"O�QqC(B������A�X"� �"O�q����V�8��B� I�Ѱ$O �,��G����O�7̝�Ԏٞ34�6�K�<@�L�-�4� �I:O"��逖6����rI���q���±$ts��M�p�S��Kt�' �qe�LYV� �&]�G�S�=���k�.��]�DE
q��%`@�#>�B���J��y`���1xM͂/�B<��S6d�0��R��:W����	�R���O.c>X�kP5��)ڠg�@�8yq�<A���`CN�.7���� :ma6���Ʌ��	9!��@�P��2�����=<b�I�t������O�a3��*?��`k��$@q�4O�S�̓�V����g�s ��],v��a`O�E��!c���GM�d��&o(�Z��:B�
	87�:�'b��!�T8ϸ�J���;s{�u��L��I�t��'��D�3oW��V/��h�< +�m ~��dڝ7� �ڕ��i���Qֈ��hO*XD��
�xDL�3��U�Q*�Њb�͸���'�l܅� Uȁ�'L��'�r�m�%�	.����Ǣ:a�܁�59����a�B��?�4Ɓ�/.��Ѝ�p��������h�2�K}~�m8�l&i����O�ptT�����$�?#<�q��62F�rE#�_���bnP~��F��?q���hO�扚{=c�F�"Syl ��P*%��C�ɢ0W����� 0A!�ǋ<d����^�����'��I�SSó�����@4B��+S��Cp`��ȟ�������Sҟ��	�|�����0��s��>s{�M��Ώ�k�ܠ1pb�(y:t�P���<���A�?�h����4~n�"&�Jg�P�Ѝ,� �B �����<!��ş,�%)�,�l�3�֖H�
Y�t$C��G{b�I�L9
 ��"�bz�p��	�{�DB�I3I�5
�$�kx~�ؗ�ҹ������'��99� ��F��h>�:�	�`P�B.~�꘸��O�19�`�O���O��C�+҈T)Z�a1AN5H�ɴm>�2.�|��s�A�!z* ҲM*�~	(!;��]�U��	�B�p4t�Ӫ8ӼD3F�3	�"u����T��#>a%�O��� �S{�586Ǝ75~B=�V��{e�˓�0?5 R�=L����?�֜3d,Hx�`�+O@uqPI�"_j\X?�J��N˓�=�%�i���'��ӹ>�V�������Ö�VP��B��Z��#�Q���7�`j���ܒ
����S���iƹ�(�y�i�U�&A
фR�+���m�x�PĮ�4(��*�'Zf=��Г=m�|p���4t����/S
��I˟���'��� I�$F-I�pq�����R�`�0�"O6Q��D+E�-���ܰ_�j�J��I5�ȟ���F$���>Ѹ��?~ʒ�P�m�Ov���O��sj��f���O����O���;�?!`I��R)�g�F�T�±�v�?��Q����Ozd���]��Xȟ�h�>�E͚�j��ka��j[����bO�k�� �`§	�`�U�'Z	z@�O}�c�@�1CJ�y�v��P��*Xyn]#�	6?IA�矄�	I�'&��בF�P�h��>���f��=+�!򄏽`�U�S�Qsܲ	˷��0�2�$��|"��򤓊G�:L� Y�"�4M)��E�f�R9y1M�6@ ���O�$�O4I���?�����ȩy�&�8��g���z(�/j����sj�ѥ�Ʀ� I�F*�E��8���K5>D,�ѓ'�$0r S�E]�<���@��ac�J*"=�������O�T�W���@��T�l���i�O�=1���Ԃ1 �{gZ���W�!��Η�$=C��U��腇Ys*�I��M����DV=���mğL���|J�	q��i���GZ����şذ� \ğ�	��p掉{b�����w6Թ��eF�s��͆2w
�#��R'#�$�Q�/�1p����`BJ�������<	�&�9�h��uw+��V��B�)�3�̙iw����O`����'�>-KS%�1 ����ē6u�(+��(D�|���G K�X��������'�O4=�'sL��j�.��T���� �0A�,O��$�O�O�@~R��nt�C��%�d�td�0<����J�/�Xt�ȯh,<���[f�O�@ِ�x���;|��4���6$"���lK+JN����~rL����|�%����c����AJi�.>��d�p�D�<��5k�O��|R�ȅT�N�ɰ��	P�>��#O
X��O?���9O�X�5*֐ez�	krl�P�5Y���^\�0��YE��O�PJ�'�6ٙB��ێ�bC�G�Zt
��'���xN�,�H!�'Rs�,P��КY��`T�A!}F��:��`Q�O�@�O@�s�>ѣ�i
����G OM��z`�L��.HK/O(Av�>��,H�(�%�~>H�Z��ߔ:����',f�N���<9�K�K~R��#�2X����Pٲ�CG�ܤO������ӀH�TH��		6����"ͪ,����~r�T����?�RX�I�44X�5��=���jF
�2uD��CҰ?!7��m�*Q�gD̹+D	Yb�D�<��eL�0+H�rc+_�r�$J0% ���IKy�'�|�P>�؛{M$TK�L w"�adΎ�Rp>����?)��(�.,�����5HI�!`�	H\|T"�"OS�Q�*�@,�<yRz�r"O|�g�ՔB�3B�\%GYp��"O�!RS	��~�[@
�2fv���"O��p�A�8K�h c�8,b�5)�"O���6�P�W
e����=S*Z�C�"O������-n�,�M>��"Ol��c���J�ny�pe�		f�W"O�\ �B	�  A���P�� �c"OP|*�V�3�(�w�A�o�<0�A"Oz������mKwdT�R�:6��������������f�ˮL8�y�Ad��q�>�KU����M����?����?)��?q��?���?Q��_JodѠf�2S��ʀiV-[���'��'n"�'�"�'�r�'dR�8[��-j�n�!�``xs���l�6M�O��$�OD�$�Ol�D�O(�$�O��$�>x�݋(˔N8ʩ�f��\�X�mZ��p�	韘��՟���ȟd�IǟH�ɪ{�x�0��]�u�@���(3ބ@�4�?���?Y��?���?���?��FHi�&Q>�����fH�	"�i�2�'u��'yr�'l��'���'�$���	D? D�G�a�f�+�#c�*�d�O��D�O���OH���O����OЁ�HO�z��H�'y��`�*LĦe��ǟ��I��������Ο��I�ĉŘI�:�so�2v�:h��qmڟ���l�	����I�X�	������I�h5���ϻk�zpx#c��qmh���4�?Q���?����?����?1��?��>7HDh��-���&+Q�i/�U���iF���i���'[B�'���'j�%���fd�Kӊ(_��9�@�7"7��Op��O���OT���OJ�D�O�����J�sӋ^�B!ڑ�c l�yn�X~R�'e�{�O��@�&�tٱ�"@�NK��-�J�oZ�f
�c�,��3�i��$�5n" ���ˍH`xiaթ��]���'^�ķ>�N~�rFG4�MC�'`�gU���*R���Vz���y��O89��4����8��d���k�*��e÷ap��D�<�H>�C�i��@y2� fX����%\,���MC�	�b��s���O}��'�<Ox�'�``�i$v�������'j�p��'�B���0�Z�O��?�(n�D	��BE~���!��)�ʕPQ�<�-O���+�g?! ��$5X�Y�1j<ψ���"b���4'R�I�'s6�7�i>��׌W�#A�-����������
˟D��(�� _ �|m�c~b0�����!�M.r�1
WMY�b�XA�hNI�'$�[�@�|"f�U�[o��Ԃ\��\�Pjy��tӊ�i���8�ӣ*:բ"L�.<Jx���]K M��O��D�OD�	E�OD�L�/2|
p[a	:T?�)��+~�d���Of�D��?�u�/�d�<᳅�v�(׊�����qQH�4��$�O&�D�O$��<ᑾi ܚ69OpUk3L�c�l)�����aZ2�'�
7�:�I2���Ѧ1��4?�ǒ�#ȡ�Th�/}��(�퇿c���ٴ�y������Wˎ&AXC�'c�Կ���;m5���t�Z4�i�3G�\)������I0�IƟ���J�Op�6���J W"�{o�� �c�O����Ot|l��+�~��I��0��4��'����4m��h\�$�b�_*^J0㑟x2�e� Tm��?E����͓.T^0/$���̔� ��8+6�0"�.���o8�XI(r�i��U�2ʓ�?���?a���Ra��C��|��n�2e�m���?I*O�`m��d�2��Iӟ���X�4�$\��C�����,kB@�����a}Ҭ`Ӕ�l����|��'���ȏ�����%���A�T�1p۴kQ�I��u7�w?�(O`���+T��a��5�:��&�d����O����O��)�ɡ<93�i�>��S&<WD0ҷo�{\��C,�R�'��6+�ɽ��d���� nI8#��yUi��w�,��%�A��MF�i>�8�f�i%���O�ٕ�+��4^���աIJȔ)d)�0�8jG$��Ms*O��d�O��d�O$�D�O��'��H��\�?dJ���	M�|ٴ������?Y���O*7~�@���n����#T?:}�i"LԦ�[ڴ`��'��$�O��U� q�61Oꘋ���];��j��<R��$���O"�𷣜+�~bP�Px�4����O��Ĉ
!3�0���0X�=��*1Ϟ�D�O|���O�˓2q����:N�R�'����4h8~i���rpa#�m��O�=�'��ir�O`��hČ�`�W@�S�t�a�'�2�)p@JU;E�i��b1�N�)�~8OI`��
�� �c
��L@D)��'�2�'���'9�>��a?���q+MB����Dk�&��ɖ�M�Z��?��%͛v���ꃄ�>�"l�ag�!s�8(FCo��oZ�ME�io���i{�$�O��� ��D�4=����F�f$�%@̬Cq�
�MC.O����O��D�O��D�O�$�0�D�g�$0�eQ| $�<1C�iC@��3�'I��'M�OK႕��5J���ǚ��&e�,B0ʓ�?a�4(�ɧ��������mB�,�4L�3�PIƕ�"����4<��#0�<�a�O ˓Ea��S�D��>:l��W��Z���Ath�ϟ��Iڟ��ʟ���{y�
q����OұbR�9�^4��ĂY(\ �D��O8�oJ������Ms�i�\��S*�b��M �JJ�!�#�]��5��7OV��D8R3u�O����u�9�ꐢa�(춡��
�B��f�'��'p�'gB�'�>�R�HU,C��[CdE�KgZ�sW�OV��O oZ�J�h��Iꟈ�4��'u�]з$Wk<�9�`�r��q�p�|��i�7-�d�zӢ�I��D��¸<��!ļ9e<c�Gh���3�Ot�>ћFP����ǟ\�	ן�R�O�!=a$��,
?���!���|�	ky"�q�~�y5n�OR�$�O��'"x�p�ԎR�H@���I�%��З'T�J�F'a�t<%��S�?�������K��łHVf<ąҴԼ������4|8�'��dJ���᠐|B�B$��t�#_���;jU+C��'jb�'�����_��Aٴj�B|��L�e�T�7c�*G?,(/��?I�l<�����L}R~��]*��<.�ؐ���
38>�����Ոߴn|�<Bش�yB�'`�QR&���?��qU���0ᇪ�e��cF��ěП��'oB�'k"�'�R�'��K�����!D��4PvΏ��>�m�gg64�'s2��4�'H�6f�(s�j�$E'�����ˆ�bs��򦍓�4f�'���O��d �:�F4O����>mz���ʋ�0�,$�O�O@쓠���?!�+��<����?y�NؿKtt�����1%k"�Y L� �?A��?������TҦaB��Xԟ����8�L�%J�D��i��\���j�s����I�|nZ��W��a�=,����E[�G���	؟(#��E�l��������'���G��z���P�W0�{v%��O�!��FB�pڀ�K�
Q(Cā&&���`�=cqI�O��\Φ]�?���K `�)aF�+��HÈ�eT�����Bg�mbӤ4n�2E��o��<���7��1�v��j�i��d�t0d 6��pPǤG�䓴�d;OT���j
�n	��b��e�W��P�4�S���?)����O��|��P
h�򣟛ZD�9�AE�>QV�i��7��t�i>e�S�?�xT�L5�![�(ڳ"Ӷ�ȔoD;B��l?��G�#��1�'��'@�	2PeɅ�E�BP�ǂ+\ƙ�I͟���ӟ8��ʟX�'`n7M��\��"� tm�BqlX�&CÑd�xD���'�87m.�ɶ���O|��O�i�g�Y�1�����JMj���/tc�5O��N�4>ځ��'ac�����w�,\���4K����1�¤dO �1��?���?A���?�����0ik��A�g\lA�@A�a�<<�$�'�'<�6M��L���O��n�N�qY��dmQ�0� ��&f��O<a�i��7m��h�qB�fӐ�����M6+�n,��!!T?�P�w�(>� ����'�5'���'�R�'���'e�-I�J��Gc@=����S�݂��'��T���4�6�@���?�����I�&sh�A;H��~���P/��Y�ɭ����ΦՀ�45҉��4�Oq��0��l#��!�+�R�x1���I:c��bE
��[��	�?���'cn�&�0���c$T\�j?$���՟���h�I�p$?Ŗ'3�6��7�0��фC �u@�
W�R�l0q���<�'�i��O�u�'M����PQ��W9�d���M*+_��&q��%�Tu�.��ޟ�Ht�ʔW���<���:\�D!�˞=]v �� ѻ�?�-Ov�D�O��d�O����O*���$�G4 A�EY�~��\Sشp3�����?�����OK�7���5É�W����@�h#��i�B��9X޴D �'��T�O��4j4&֛�1O�$ �ř�M7ʔ�W��s�^�e�O��Jr#��~b�|�W���	ٟ����9�0�6I�IS<A�V⟄�Iڟ��Xy��i�ju��D�O���OΠZdI��5/�Mr��K�rn�hۅ�9�ɗ��D�Ħ-�ܴ/��'h8eA��.}�m��'�V���:W�'&�^�lC���i�Z˓��⠬��ϓb�,�@G�1W�ɑeBZI�J)�	ǟ|�	ӟH��x�O��D�$ꐙ�BG0W(�U/m�"�~Ӡ	�wb�<״i��O���9���L�=$�hp,{�^����͒ߴm����A���<O$��\�B������\�����9X����[{҉ R�$�d�<!��?����?���?	�F��5��ݻB���'�4�3)�3��O�8��ݟT�	؟@��N�t�']0��%L� ��m��F6���3�>���i!h�D:�4�V�����|� ���\@�s�� Lh��Xq������5�<�Wc�1y�(�$������\ L౎P+j�v1��DR�$�v���O����O����O�ʓaq���	Q�Re�h�zBg��T(�3�L(�jg���|��OV�lڜ�?��A?��7ͅ��m:���1G�y3U��æu��?��P5G�`�������&�ݧL���r/ޟ^Bx��g�>Kf8���O��d�On�d�O���<§zSj�1#�Ȟ^y8\�5K!r�T��ڟ��I.�M#!b�������<�c@Xb�i3AS�1z��k����ēa�F�m�����	~��7-u�$�ɜ:>p����y�r�z���C��!�w�°*��/|�Ipy�'/��'�b�]�nG�5)䄃1.l���n��0�b�'�0�M�׬7�?����?	����$��J��4ae,_f�@�!���D�W}�c�P�m�%���|���l�����f5a6n�S`H���l�5���>�N$jbCF6������Hr����O�����(����EՔ7���m�O���O����O&����^�����^��온|�����M
�1�>8�A�'�r�oӾ�D��OLtl�ox�yj5Ϝ�!�\p�Q�ҶV�ĉ����M����M3�O4��c�RVi2z���SL�� L��NW\4� �Y�d�'+B�'��'"�'��S�?����8��DX�@�@lz�����'���'p�T>%�	=�MÛwf�sG�M�  ���MкU��in�6m@B��?-��?�KM�ߦ��w[d��䂿
x-I���	�����#M��K���OV��J>Y(O���`"�2&%�&�A��D�!n�h!"��O����OzpBT��k�tQ2�Ô��� `�%������Rܦi��4R�'��� ���%UFb +�{�FԸR�'t!� &���Fb2��I�?����'5���Oh U�0�-c�l���%LR�����Iȟ��I_�OF�d� �X�D�ȨP蹛PJLhZ�MtH(�?9��+����$�^�q��J+|�j(�&O�A_P�{� �O,�nZ��M��i�6ݑa�i)��Q�Ē�ҟ�Q@V�� ;$ ̪��_�$U�]8��:���<���?Q��?Q���?�h�2]ZD��n=-!d*�$������(��P�x��� '?�	#wP���CM!��C��)�OH�d�O�)$��Sݟ���.Y<�`��_!=�ЛF� �FHB�� J���=k.Ot4b�]��~B�|�^��*��x�Гf�V�V�����@����������۟d�ITy� rӾIR��O� �`i���j#�Ӈ}f�[�hڹ�?IB�ii�O���'���'����O# ;��@-���(J�GͨVT0���i'��OԨ9��L���Y���߼[􊃣:7`��ƭ�6X.��gύݟ<�I˟�Iȟh�	�E�ĩ�R�e3Y:3g���*�>�?��?Y��iJ�i�_&��'T�7-)��]"�|���� ,�X���?N�$�X��؟��<x�Ym��<)�O3�� ��T�d��y�� C%I7l�y�D�J�D��G�Idy��'�b�'�N�o��+C�%T�r��C؇H��'��	��M���7�?q��?�ɟD}J�숻mk� kG0��ɰBQ�tI�O6po%�?)J<�'��W�.?6ty{'L�����C�� �@�"���(\q܈;*O
�)��?	#�!���/_�|*��(�P�W�.m����O���O��$?��<�6�i�� �}r���}Ykũ�T~���6'��'�$7��OēO.u�'�:7͑;CyVL���Z\� ��i��3`�oښ�M�3m@)�M{�'4�"�����SN;�ɊU����a.s�6����39~ ��Zy2�'�2�'A��'��?Q����
2��Y�S�ѯ\�j��&JIʦ�Q�eT��(��%?!�ɠ�M+�'T�9�h?Y��c/A�{��#r�i@��"��\�	������mӚ�	������I�xs.��1eǐ@��	�I-�ͩ��'\v($�ܕ'��'�h��׮A]���e�-��b��'���'v�^�8*ܴS�~A���?�P��ܲd��&�����),�p��`�>�B�i��D6���*(���6E@ ,�NA�/ٖe�.�d�O���I�+~��l!��<��3���d�"�yr�]-kn�z�� �s�l��'��?��?����?����a�� 2��4|��	R��g��xk��O��lZ�
xHI�'mH6m*���?M��DН<�&�gd�%-�D����ϟ\�۴!⛆
k��k!�t�b�şH�@T
z�TD�7,+�a�7O˕�4
7��
)@�&� �'�axrO�����:b�I�d��b:�'t�7Mϖ3�@�D�O|�$+�S !�nm��@�c-�-�$H�X�h�O�o�:�MS��x�O����Ov�]�/ZS�Pyb�2x-\雲!5p-�V)�<A�
� ��	`�@yHZ�GÌ���%U?j0Lt[5	$+]R�'D��'�b�'��	��M����y��Y#.��� f�~�����[)�?9ýi�O�L�'�j7����Y���@1"1���j��-[�)C��X��� ����̓�?��
+�p��]���,�$4&L#���>>}�q��	I�W)�d�OH��O��d�Or�$0§O|���7N�(#6�T�U�Ӛ!���	̟���,�M[!����RҦ��<wњ/�"��&B�xx��1�1�ēV6���g������v�6Md���0p?��J��{���C7o\*U�V�Hlʄ~�2��m��Eyb�'���'&Z*`.:� �JC%3D:��ğ���Ty�Jc�>(ITH�O����O�'���8�O7D�y�&ʛ���'�Fʓ�?������?��e��@fͰ(�QPd�^;�����N�*,pYqBWyR�O/2��	
y�'+Z���¬G3]8�c���|��'��'��'��O
�	7�Mӄ�U�L��	 �W$}T,"�ki*��(O�mmZ{��xT����M�B��o� �c�oo8�k��C#�fHp�d�� �oӈ���lTٖ��4�^ay���%6�s�"�,b��K�+�2S���I��<��ݟ|��ɟ�OS����Er>`�B)$�����iL��` �'��'�O��gu� ��!EЬ��$N�21x��Ešm3$��ݦ�RN>���?��S�a�*,n�<��ώ�V�L���%82@���?AՋ^,S��I@�Iiy�'-2k0m�	��E�z�V �Î�$W��'{�'�剼�M���=�?���?ц73d<���ӶqJu
�D̈��'����?���p�'f��/xb-�F�ʈfVV�jP�վrD��'l��i���=��f��<q�'���I�<�2�ȵX&}H+H>!`x�OD��0�	ʟ��I�G��=O��!���"%A�#S�4����'F�7M@=	)x�$�O�umP�Ӽ�L%Tu Y�*S3�p��cZ=�?A���?q�i��T�i��b>��c�M����ӧ`��wO�89���*D��S!�'��	ȟ�����<�Iӟ\��5ym���e�پM��<���[es.i�'�L7�ފ���OF�D>���O2i����:6���+n�E�4�FE}��'��:�4�����*t�ŸT���,[�;֤���eT\��$R��i�˓,��RW��:�?AN>A��|J��j=�4���?"B�A���?q��?q��\.�3���$�˦���M��𛡉*��e��.���9ԍJޟ��	@��ޟ��' �6�D�?���%UZX0���
l0&݋�� �`���F`|�<�I������J��!0��wy��Ogg��;0�!3GL�a�4q���|g��'gr�'k��'.����nu"M�}Lj!����%[�V�D�O��dR��en�KyBd`�4c�4���ڸY2��QRݏH�T�8E S�	��M;Ӳi+�T-��f6O���O]��}`�M,@P��A$@�������V��*�5���O�i�2�'�r�'_�`�g:K�(ɂo�>4V����'�W�l�ش.�ഺ���?�����iʰs�^ ��Ɉ�~e�<����V�����O�ʓZR�FJ������)�,P��.�Y��A�E,��v��	���L�Bu(i�\�Bʓ����Ox�CK>�5,�)sr���ܷ0Qڱ����*�?A��?���?aM~j*O�o�2H5�wi��{��r���\k<���T⟀�ɤ�MK�Rʹ>���i�P���#�;����J�%�l�Je��n3ApJ!l�<i��`�1t��:,�*Ox��$�93�`1�@�%A��u�E/�OJ˓�?a��?����?����	�3ڬl�b��'_;$��:6��X�D�O2�$'�	�OH�l��<�a�I�,ZHSĎD�\h��Eh��?�����?���?�X�H7i�$C#O�![,$���QFJ�8'���$2͂�iR���]�	Tyb�'�B�6M��s!D�1,؀�g�-w"�'
R�'f�I�M32 ��?��?��������P�/��P���+��'k��k�����*X$��(#��\�Ĕ1�*X9�����ky�Ę`|�Cee*��Oa�9�I*���6cbP=�ǇN#�:��1��f�b�'D��'���<� ��S1fF�/}����}�D��'E6��'m�v���OBYmS���b��#7�B��c�[s��� LO��?q���?Y%�iKhdZ&�i��Dx>�YA@���dnE��]8s.R���P;���

��'����D�������Ο �ɣj;D�9^�QwJ���=nw��'�<7�J-U���?YL~�;8���2C��Τq��[�p�N�'\7͕+�Or�'���'r�2!�W�;%U��흓G�L;�&�M�&P�<Q�N۴nm���R�wy�$�<���yUDP-26"���Ӱ,F��'�'t�'���M����?!�oΐՀ�A�#{�>�V�?9�i��Obx�'v��'���D�20��5�3O�2P�8-
1�G'�����iL�$�O&�H�DY����[�D����6��?�t�G��B��������ޟ����l�	���D�4�^�]�sQ��t�KfG�9�?���?!V�i�$$0��'�Ayӎc���g��P�0��#���q4�ZH�	���I�?�[ڒͦ�ϓ��B�=~�ڕ3â��a2F�x���v6�y 3	��(&���'���'�b�'1� ��-S�q�zp�t)ν� 9s�'�r]��kݴ&�p��?�������#7>~�;D�1}��Y�,8R剰��d�Od���o�i>��	Y@:�I򍌣+wd�9��1!��Q�E�Ә|�2�lZ��������[�'d�'z4��t2�Y���R��Q�'���'q"�'-�OQ剀�M�c�f��88BI�W�]���Z#y��@���?���i2�|"
�>�#�iH�!bvG�56;0Q�ȅ6fi,!�!H|�dLm�>9�l��<���8S<�)��럾1)O��D��J��-�P�^�ؕ��Oh��?9���?)��?9����)�;��!y�$X�1U�Qď�~+x7�С	n����O���!�9O��m�<�t��E�F,��eΥa��xh�MP����I�ē�?����e���M��'��@@�D(7+�hJ�'�#?E�I�V�'J�s��g?aH>�)O��O��[!H<ꄸ��A�P0����O*�$�O����<���iq�0���'_��'H���ڙ^m�ۤC��Z���Ї�d_y}��'��c)��2mq���!�F6I�a�V�Y�<���$�O�TA�D�j��6�Jy��O A���yҬQ&�x)��ѱ�F)ó�ɗ�?	���?1��?����n��;RI҉+<Lpv��p� 5)$$�Obil�;�lQ��䟬�ߴ��']��+�Rt�T#�\�Ң�#<"�'��aӮ���q�(�I�|.Th�P�O�J=C��M9n�����8=��p7�|�X�H��矴����T�IП<�V�JƂ���B���UhŦ�Cy��a�x��/�O��OX�I�|j�10�(���5I{������Q��)��S���I̟�BO<�'�?!�'z����ӡ�'��1��s����	���M+bP����鍧OE��)�d�<q��ɠ-�\h NS3wD�@�5c֣�?i��?���?�����_ަ9�'ˑ������ֹ>N�hsN�,m7&�*�J���`�۴��'��ʓ�?!�4nRPB��2`Gģ�1�fBx�x��4�y��'�L�cQ�ar*O.��{ޑ�`B�j�r���N�D�)��b�O$���O����O����O*"|T-�@ld���ي~�B���I�P�I�� �4|b%i���?y��i1Ȏ����IG�d7,�"-A|�`��<�d�O��������/~Ӡ�I�|2B�F��A*� g2�i���2,�x�r��O>�Od��?Y���?��^�^(���t���%,α�.ը���?).OhLnZ�Lt�������IG�TN�U�|HN�Y��za���Ďc}��',��"�4�T����E*2#�)���\OR( ��E�%��uq�4��?�8��O��O^��!��Rِus󏎢tA��� �Oj�$�O��$�O`���ʓٛf�ּQu�@�sL�J6t|��КR˪)�'���f�r���)O����27Z�JrnK^4�zTH�P��7�O������Γ�?��A^4��ף��D�bLޅy��ȩ! ��O:;�D�<y��?���?����?aʟh�&�&p̵���Z�sq� q'aӄQ�ń�O���O������ݦa͓@NT�E쀗}X�TC�@Ö{�� �4<���E?�d������p��A|���	.=����j@a��)�y�4��	>0f�O��O��?���g�Z���&�*�(�j�D��`�	��?���?�(O:Tm�aOV=��ş��ɌB�uc(��2�41y��j�-�?�]�t��ܟ8qI<��)U�,!�\� Q>g�y%���?����Q�I]��M;rV�����O���e�DC% <��Ё�Mr$d���O��$�O,���O4�}2�'�$z"�L	HtH�� ��
��3/��юI��I��M���O`�05	�6c���Ю�_K�<�g�'�R7M�Ц�bشu�b�j۴�y2�'��%E�R��J�?g�2Es�!�s�h��e������O��D�O����O��D� e�|3���1D�@k��I���J��(�Z?��͟��B���&�Q`�F�5X̌���^�%��	;�M�׼i9�O�����i�*`y[�	��f�hR��"����r�^�'C <�e?IJ>�*O����@��
���eG!H�D�i�OD���OJ���O��D�<Q��i�fS��d��O�܂�N�{�x`d
G���I��Mk���>�ոi�7L͟���.ȷ'w�3s�
>)!�T�ͱs��7�h��	�
�~�7՟P˓�Қw���(�N�{بQ�G�Uy�ň��?	���?���?����� .��c����	��q8�:vS�T����M�����?���&�dݓcc�H$ܐ(�^�x�a�>V,�OH�n��Ms��5v�,��4�y��'*�:�煞)xx��u���!�� �R�Ј)X���	\n�'��۟��	ퟀ�I�vXH�36���Z��*ᢃ
MP�����P�'N7�C������O��%����*ҘZ�i��k�F|�PP�'����?���T+���T�'�N���AĨA����-�h�m�&t���p��F"�M2Q���%]3�D+��Ҧ-�Y��;X��)W�J��d�O����O6�d8���<ag�i����4Ң��)��n����.�Q}�'��7M0�ɤ��$�O���æ1 ��$�Z#�,���'�OKh�BC�b�V���|Ҕ$F7��ɻ<�P�֌���0��8s��h�g-�?�(O���O��$�O����OZ�'x���;x:Qâ�Yy���4Cc�}���?�����O��D�O\���*����ԛ�����
2՘tlZ�?i�O~����v�	�^���r���I�L*!�� ��5���Z'a�X��	#z�\(`�'��Q'�L�'���'��I:D��?b2faA������s�'�Z*N�����dЦ͙&���`�	ߟ���܂U�0�i�,	-N�2�*pm�~��ퟬ�'�R7��ßx�'�]M�LŢ�B8)�t}��j��+�r�'d����?,m� Y�T��1�b��<	�"��xX�x�d#8t�9�b��͟��I��I՟�E��2O��J��A0�F�	P`�)B��'%$6M��%'��
���D�^�㲅�4�hj���d�ޥ[u��O����O��m�}]* oZ~���c�Թ�'þ�{���d���2H#=A:�I>�*OD���O����O��$�O�u�V�d`6�{Sc
(E�����<��i�i���' �'��y��� v��©ƎAB��m�(\���^7�ft��+��)&j��qXCÌc����ĠA�-�e2$ g�ʓ1&Ц-�O�	�H>�.O4�Y ��0?�Ȁ �W�	"k�O���O@���O.�$�<yD�i��}�5�'BD�,ݔ[��8� 烒2��xٓ�'��7m9�	���D�O �d�����p��֤�d��]q�Y�M�%J7-0?)�Y�l:��H�Sü�"Ξ8mG����9\>�J�I���Iܟ��I������hD�d� @�z�g�3a������Ǎ�?����?A��i�����^��۴��'6�:F� l�.f�]��2���x"�'�"�O� �iu�dv>!�&ʛ�)��р$Ѐ5j���Ѯ�; %t��'��'��I���I��	�l!X����8n	p�c��W�����4�'�$7L-��$�Ox�$2:Pą�+G�)�s�kת�s�h
hy�#�>)��i�6��U�i>u�L��q�@�,2�Y�J:��d�$��V�x�n�����޴b�'j�'j��� \-$ q[SH�Nr� '�'*��'Mr�'m�Oi��M�F�g �͠�̆���qᎭ5�j�[���?Q �i1�Oxt�'��7m;�*=q��]�X@���.g,�m�"�Ms/�M�'�2�	�������������@�(�a�m����Q�l���<����?)���?���?1̟��`�	�L�Ip�M&=�¼:�)|�Ľ�C�O����Of��|��Wn�f;��Y#�E`�f��g��D<�}�4�lZ+�����'��M�M3�'f| %��0�^8���ݣB�8��W�'��xC��џ(*$�|[��'��GN��8Q��C�K9�����Y��e�T��T��Ꞔc!�_!f��A)�egnhR!�]�V��I��M��iW�O
!"�I��G�y�7�΍L�T�0��OL�D�73�U�bx���'��$�V?��'�ڠ�q���S%:�'�#QXz��
�'B������Yx�@V)żxZja��'�vHS�2�'(�6&���?� ��ӄU��f(.^�X��f�<QݴB����w�(K��x�Z�I��굄U�j�i�)mhPc�֋W	v�r�-P�<�O~ʓ�?����?����?���*�Q�&؍Ej�H��80bMB(OH]m/��I��	c�s�T���S�u�F-��Ѐ4<��@��Y���d����(&��S�?���&V����N@'hT�xx�T��X��E����bT�'�z�`�֟����|RS�t*�]#�2H�ɽ=�PQ��+ǟ|�	ӟ����@�	qyB�hӜ�Ѕ��O�q���T�E'�Ӏ>
vI���O2�ma��Wu���M�1�iG����b
���Q��C��%]ߖ���l���?A��������}y��O
�N *&�(���0���:U�X?]�r�'��'�R�'t�S�d$�ǘ�*��s���[dʓ�?��i~@0�b�'0�u��b�d��+�<���#�A�jY,L�Q��V�ɳ�M��i]�dMC�u�=O��dC�-� �S�H	8t��ar�*,tr���»�?�C2���<���?���?�"NZ�R7������ ��`���?������� &Y�<��ȟ��O�h�Ap��u:���ьy�PhS(O�u�'S7MU�)0N<�'��B`H4Q�d��H�5&�5�Q�ԁdE�a��"?�ޔ#(O��	D-�?QS�)���6O9 � �"J�E�l;�(�0���O����Oh�d$��<a`�id0�z�E��9�`�0rțK��q;�! X剮�Mˍ�Ȼ>���i�R%3�O!;f�%p�I_�t�Ja��auӖ�m�`,m��<���k~��C�����S/O���G�].>�����OҲL�$iX"��O�˓�?A��?����?I���� ���@�V0]��-�PGߣL��P,oӰU÷K�O����O̓���$S����d�he��˚A�:qy��&`�YS��?	L>���?����e�2(mZ�<ɒ��ك���'�p�&/Q��?iA���&�����䓤�d�Od���J��}`���f2�BɫN��d�O@���O��Z"��bJ�:��'���\V{� ��t4�� ���?#��O��'���'��'��)��匨y��G���l�0��.O�usL@��X��3��=�?���z������ȩ�0eW�3���D�O`���O�d�O��}��'�>���L@9��!ڇ�2l&�L0�*����D���'ۮ7*�I�?A1�!��{��R�:7�J��ʞ���+شy_��m� �p1�a�T�I���c���;��T!�*g6|iɂ(��q�lT(^",'�Е'���'"r�'���'L�K $�7! 	�#g���Z��V[�8��4{��8(���?I���'�?���0x\8��KL��1��C�O����nZ!���?���?Y�j�^I�}�B �&ss`U�T_�5`"n������J�!�'��' ��'�ܨ�&(ǃ$�U�EŶ���	�����������$�'ܸ6��2u��Q<%��B��܅FP����g��b�����즑�?Q�[���	������U��Ώ(��,�`E����$h�EЦ5͓�?�#~��Ly2�O���ܶ&��b�H�;��\Ӵ�ÇK7��'J�'�b�'���#tQD��2i�1!���
U${rʓ�?��i�����O��9��NT�qĦH��a�����]�:�'��$sӖ�oZ�?��������?�p�	6��`�$d�'(r��ӂ+� ����?�H>���|���?1��?)��X%ZvU��nˁr��(""�7�?���D�Ǧy�Ƌ2?�������bt�ɿ c>@*� ҹ!����(O
ʓ����z�
��'���?�����A�[��,L�8�1Sf�lH���MΦ�/O$�I߇�~�|�O�&UNL3�	���p�g���[�"�'F��'�2�'ذ��H�:j��	��M#�F�+`�����@A�L2�4@Ǐ�b��"���?������?�,O��n�T�ڵg�<s֡��`":#2ABݴI㛖��%I��=O~�d�8�M;wa��?�'���ԃۣ|���8�U�j��ؚ'8�	۟4���|�I��,��T�D˨J�~9怅+A��bG_�B���O__#�M��'H��OUr �u�'\�'�󄔈`(Q�!'�r�D��J7-R����OV����|��韮���q��i��P�����X����Ĳ;2@�a�i�� q�V�~b�|2[�����,�����eM���ŎQ}��Y7� ��\�	˟���Iy��~����B�OJ�$�O* *Uk_+J�YkDH�+T�H���:����dئy�޴��'�E�֤�7Wx�:e�ߞH�L�"@\�H����X�Ll������I�<���	q~�x	E��xn �3
���ҟ\�	ş�F��:OhaILT/,��t��#��i���'�>7�K�H��D�O��n�{���r��\�KJ�=�C��|R�ɘ�T��?���i�p6m�Ԧ5{��KЦI�'��L�тM�?��G^�BԺ��&<��;Eᄈr��'�����IݟX�����M8M"�lX�G��u ҂�v(�'&d7��((���?!��TJL<.	�	%M�j�b��{ĲIc�V�H�	��+N>%?�	��-Bڝ��朝S��(�� �0p���r��{y�R�$�Ƶ��o��'���)�uf�.s�P�+��ΏL0�8 ��'QB�'R��'p�T��Y�4]����$�H�e�+E�$XCRjA�5�L���^�6��BT}��'��/�O�8"�-# ���D��%�t]��D�I�6����5)Խ<���<�I� G�J%P�Ɣ�J��aJ�()���M����x�	͵B��ȁ�!V8�����%[!�0?)��P�Nm�	bШ w2����
 ���*$�)�\֢F#����Q(ȥX֔A�Q�Ůk9Bd�@�
����? ��<{�H�(�����X�U�t�U�]����l�DhD�]�T�25�dK�4�`=�Pȗ�NM	(�힨s�@��#��a�"�gD.x�<R�HG�.垲8XiP�U#U���'���bR��b[���{�mW+a��up��یsh��j�'�r^�d�	ߟ`�����'����J�4�2�/��NV�8�h�H%��Q���O����O2����9j}h�� ��)�,�	&Θ�c	�@`R��v���Ab\,x�@l{6ON�$�O��4�P6M�5�V�c�o���岡n[�w4���l�Ioy��'�`��t�i�l$)�F0�B4�)V��}k�'�2�'�L���'��/x0��'��$�Mx2~�ˑ�0,6�8�l��;P�0dT�1�"��'�2�'Q�O-�ğ�'�u1��=\TE�S�ޤ-0Hr�'k"� M��Q���I�?�O�	�s�]�77j�J`G_�D����V,�����LI�wy���Iןh2�@B�dJh��䟰����@�ѧ��<i<�R�FH�t���@����3w���P��ٟH�����'2�i�zl�P���	Gle���6����,�<q��X�&E|2�'�&���4@�b��Ur�!�#i��kҠ�d�Z֖AC4��$<��$�O�) �Pr�1�19O�6�
;!�{�M�S�d%�<��4�I|y��'�B�'�BT�0�ɜe�du:�*ǟJ0Й!g�&6��t�)��?I��?���\��Ⱥ#�8@8V�6I�:!N�8�j�/�@�s��?i0k��o�,��6�]�<���?i��|zݴj�f�ym�Z��)��A\�I���'�r�'������ �k)�����E��N��աO�:��E������I��$
p����sP�,����I�?ي���}�� ��Qn��&gP1 &���P2�AR�4�	矀��ʟ��ҟ4�I����'�,��X�C�
��B��56M2��'>�!�&�Y���	�?�Oh+��H��ҕ1d��2����CN�%�P���_m\���a"��y�������5q�f��
�9W@I�1�d)k&�R;p��I�ޖ`�ة{�Ƙ�P���W�B�)ɜ���[�^Y�%z4��4o�|H�>y�.ñ�h���>�$py���P��e�d�J� �!qY����8���� �"�T��R�k�F�����<Z��MYc!/Z�:�v�G�s�xuJڑ;
j�%,Q�y�$�:pČ*N����# %F�J�8��@�[��zQ)\�R�b�ؑ�Ҫ
5s�LA�)ȡ��m��P�������&��'�(P(`a�-HO$��B�		O���s�'�d�`���S�0⡏!�D��,Y�!p�Q�O���M���?��Z�(͑g�x��'4"=ON5xAh�%�L�1b פq+�Ds��%:\h�<��?���B�e���ؒ�A�.N&J�$����?�҅R:�'���'T�'�����J�'�* Z6�[3L����\���À1�͟(�Iܟ4�'�q��g�9�(��DK=Q��1��X�.��O��D�O.�O�ʓ>2�*���ֺV�TNt !���>]�1O$���O��D�<і X'g����r
,J1 $%E>�l�2
�I˟(�	Q�	Ky"L6�~ X�r����L�"!)��A�����OX�d�O�u���s��DP�P��kRсP�L��B�G
���'�'��ɦ?f����&���G��(C���)gl�O���O:˓B_���V����'u����4 {,;�m^�+;�(���*X�W��'P� 0ɟ�i>�!��$b�� c����b�*x�G�'��cy�}�ش��i�OL��REygX.��X ����XC%ɓ��?�*O�YC�)�S�
pʽ��Y�oX~�$"���Vt�$Xn� �	ٟ����ē�?)�Y*lAn-�FE�iI��rq)�2�?A�'�g�����Q��;��4_�\�T(� ���mZןD�I۟�2 ���')21O4�)E	����B�*�`k�:��'�
$ӎyr�'�"�'�T��e�Ҟ3CNeʤJӞU9=�6�'�,2Lb2O�d�O��O�[�`_�����?�4p��/�<&@�m��?���?�(O�%%�8�*l�G
�:0���>tS�&�|��՟�$�x�'�t:V�E�(��cX�r֍p&%�ۘ'B��'��X���0�.���N�%$$*�˙� �����Ο��'C�|r�'B��783ri	�X�:%��)�"$+�v��#(OZ���Oj���<i�b�	fc�S��� D�E�.dڑ�v�afş$��n�Iş �Ʉt}0��<�ꎱ�z�cVΌ�(!�Eϟp�I����']�ゥ~J���?i�'s�"�7.B(+N��`��
�F�AM>i���?����?Y�O;��唁��@$M)D�Yh������4� mZ�T�	̟����B#,�q���E�0�JF9q���O��D�*���|jфT�'#ft���M"G:��@��ԟD�5BF�MC��?����*6U���'�T�f)�/Pc��b&B$f{f���'�izv��2�S��p3F�گ8kJ- �k�':(&88d.���M����?��o}��b\�(�'_7O ,(��Ԃ}^b��Ƌ@���w��Y�ĒO�d�O���_�/dF��D)?p���F��j�D�O�}�gZ}S���	n��(O�j��$�G�Q�Ʃ�
%�'*�*�y��'G2�'y�I>Urb@��P�|_� p�����؃"�����<����䓷?��xM�D��C'1vh�0-R�7�sK� �䓯?���?+O~�#0O�?��tl (�Ɛ��%�&Pz�Q���O��?)N>���?����G?�f�\0FJ��[�c�=��Kky"�'."�'�剬��#��P���>'�4�ié!
��y"�1ma����Op�O����ONi�G?�	��-�	3���ZSO�&�����O$�ĸ<���$vG������?�X����2[ �z�%��g�aӵoAn��ԟd�	$���?ѝO׌����+'0�/N56�R�Y���Ԃ8Ԏn�ߟ���ӟ��Ӄ��dL�t�n	iV�ݜ���B�Y����O��d�%.��>�d;�ӁJ�HB`��z������h���Ӏ��l������ߟ������|*�a�u��͐�n*d��-��.���?I��?���S��'z�j��*|$x�$��� � �e�.%p6�O��d�ON 㴄�N�i>����<�r�^ D�"1���H"�)��I����Is�I�� �'��'��e�Ыg�؞o�Ȩc�XLl������b�6���|����D�O�8�끝<P-��E�\F��P�3���OT��?����?Y)On��鞍!,,�eK@G�DR�-m�>�$���	ɟp$�ԕ'����!t%�a1t���`�����'��|b�'���ЬF�|���_p�$!���<��H�A�Jϟ(�I֟��?�����D�
��k�J�_0=�U뒂`{�8rf9�$�O�ʓ�?��-��)�O��w��2Q^��"�3��b�C�O�L�Iay�ƾ��5�q����"�ʬ鳠J}�`���Of���<IP��OT7�$�����u��Y=:(TX�|�T��3ŭ���$?u�g�? ���A�P�Kv&�)��z���0�Y�����J(������Iߟh��kyB�Ջ�iՈ��-fqAc��=�2�'�R��(�6�*�y��d��vvBh01�.�3�� �?�V���i����'���'���c<�4�ޕ�f�S�PAS Dd������OXt��O�D�<M~�'�T��s�N34I����jM":H�YS6�'�2�'����e��)��O� jW�ޡHj�q3�	��8ź�����'�.��g����'�R�'��XƔq� 1+�g�Sr���'ari�:B��O���O(�O�P��6(� �P�x���@μ<��Q9�?I>y�����O��Hv��#uX8Jtf�  Pq�GO�B68˓�?�����'�"�'V␙�i�,3��	Xi'��:�O��H����$3?I���?�����[;�I�SD!��
�-�~��PZΑ�ty���<�����$�O��O���3O�!@0m 1M*���
U�%a�ą�O���O(�$�O�˓Pv��S?��;%z�b@�߬P�n(���4����󟀖's2�'���-�y�'��C�)�E�#h�]qB ��S��B�'�W���WIF0��i�O����r�a��Ha.l2d���q���Z�`�<���?��K�����9O�擉� a��Ā��VX��fR�cXz�$�<e� N�F�'�r�'r����>���	 p1T12h��~�V��3�؅�?	��?���<)*Or��?�8���"EK�d(�X A럊�z��fQ�n�П��	ϟ �ӟ���<	�Z5T:�KUo�+�����ų�?��
R�<Q)OV�d5�ڟ|Z��$�:W�F)A�i�,��M����?!�H��Z���'�=OrTi��^�/CJ�уG�*�@���'O�'�ѹ���'��?������U_���#C�ۙK��[��'.rB��2|������O�ʓ�y�bF70w���U�)o���V����$��D�O��$�O4���O��h}ȱ�3��~��l@ ���\6h$kЍU;D��	@y��'��I����I۟��AiψkohU�r�Z�7��t:��A%�8�	tyB�'*��'��I�3�J��$�P�	��E�2�D��@H
��U�I_y�':�	ߟ`�I�� #�C����M_"X��F1$ܒEYAśПP��ğ������'�l���b�~Z�wZZ}�1�V�kZE����27q��S��?!.O��d�O���G1 K�d�|�bkL�Y��8�ף�a��;�K�:�?����?y(O>XXas�t�'F��O�X8)��D�?QzY
$��q@��1Z�@������L/����Dt>iP!/ߍ��J���9[,��se�O����h%�i�2�'yb�OU��|��E��h�K��Y�F����8���?����,�͓����Oh�@P�­#L�"��	a`����@u��T�i��'{���듉�F�Q���Sǅ�	(�5��'aux�D�q�d?�$1�S�����(>���E��ip��0uN��M����?I��w^��Q���'��8O��#��0O'l�xf͏�:�P��a�'KbR�P�V�]�������ȟ4�`��Ӵ�e�
t��B׃W֟��I�.2���O���?�-O��]�P���c@�_RyB1ED&��D�O���e5O����O��D�O��d�<�� ��왐�[�A#�y��'\�r� ��%[� �'��Z�$�Iş�	���9q�"�l(�F�?+*ma�I~�8�	��	ݟ���y�Ğ�G�����v��icHޛp	�<��O
�_��X���	{y��'���'`�Ѫ�'�L9h�$�1O�Cde���,�BG_�\�	ޟ�I}yR�F�D���'�?Y"gПj bL�ʬ�01*���?������O����O:@bV>O��n����I��<�$�H$�[3 ��I�T�IMyҦ�&:^:맞?a���2U��S҄����T�0�BG9����OF���OH��e<O��$�<y�O�I�*��	.)��@E�/*����d�+1�29l��	,�S���l!Ҏ�]� 	n�WĴ�����O��$�O>,s�;O���<���t%����hQ�U�B`.8���-�?ѥav���'���'j�d��>�/O�
7 H�s����Do|Ż��O���5Ox���<���'x {��>���C���,n�� ��ob�x���O���1${@�'��ßT̓���P�--\�0���
ٔ �IɟԖ'��}����T�'�B�'#2iZq��V����蕟Ʈ��v�'�aE=hpX���$�O���yg�%w�DE aJ#mR���L����dXi�$�O ���O��d�Op�/��HȀ,�8&b6�hb-�L栴[Q%Ƅp��IQy��'��	џd��ҟpȅo_�Q�#�1P���s�A��<�	���I�(�	ğt�'O,�{�䟊Tj�3��yh��>zK, @�'��I�`�'���'�R�[�y��?G�� �����倐4D�Iڟ8��ߟ�'������~j�#��(�4f[�S\�	��NBU������?�-OV���O��D�/~h�$5?���]�T���#W:8N���d�����	ҟ��'�>�a�K�~���?��� ����"O	n+P1�֧,.)V�3(O����O����O���;��`>ё����1i�&R���t��O��m�L�i���'���O[��xMD�I�.>V�l9CL� }����?i�C)�L�')�IX�'	)��0��r.<�$�ԍߤm�ɬ1X��Qٴ�?���?�'B)�O�(mQ12| i@o��t8R��E�O�5��O��O�?]��w�? 
���Ś�l��|C���.0 X��`Ӏ�$�O��ڔF�D�>����y�CW�����U8��$��/��?aM>�t�� �䧺?���?ye�2TbdPr�Y1n���ĉ�1�?�M�#��xR�'�RS���;X�6��W��0IҐ8���&z�)�'�.up�'��Iߟ�����x�'��#���8�҈�V�A^��H�MΨB��O��O��O�$�O.�Rtog�>u�1�E!j����!��(H�$�d�<I��?����;�����+a6ᨕ���m<%H�/϶�E�|��'h�'���'���'����&��+8D4�V$�r5:���_���Ißt��y���i���e�UF� Y,�Z�(�	WY� �O6��0��O4�d��k�0��0?�עÕj���+��7����������|�'a����:�I�Ob���/���
�kދ"�B���@�=�<�O@���OX9I^��|�'xA<�0�U�-�Z= ��������'�>Hi�e���'�?Q��{/�8A}>`�D�V$C��٠�#\�T���Ol�˿p�L�|BV�ʳ9����"׫25�k1�Bß�ap��M���?I����x��'��ʅ�@�?�IA@�'^�#1�'64(�'��'��J�d�]T�@�F�F���6�B&,�>]m������՟�������?����y�%Bt�q���"f�laq��4�?iI>DǇ��䧡?����?Iq����x
�e��Zh������)�?9��4t�h��x"�'|2sv���	�eDfp"�ߨ�剎5��IKyR�'2�',�ɾ);��d��N����+�C 4� �Y��'�|��'�RyGH��� \0`Ijr��f�$�e�'��	̟��	ן��'� �i�'�減��>�.������{�&x�TQ����ʟ@&����ʟ`���w���mO�@Ĭ]C�/0V^���&^Iy"�'���'$��)W�2QK|B���X�K�	Cj�:2%��%j��D.ړ�?������?1�O�QHBjֈQ�qA�dZ�s���B�'���'J� uI�0�M|���ygG�5@`u��D=h�@�&A6��'i�D�b��|�Old�m�D(�ġ4)�:9@�}�����DZ%n�bm�E���'����<y���X��u���M��$�� LCy��'���j!�';ɧ�O���⋍�6���9Ev4����!D,9���?y���?���?!����I@%f�p��Bt�
�Ď�H�j�D��Љ�p����dJ�;�B��Fk�2#�lR����Mc��?A�'����x�O�2�'M�Yv�H3HZ��
��½" z1
 ���v1O����O\���zk�TR[�L�j�)"@\uxa�'I��W� ��l���'��'M���g���Wd�L;č�Қ|�����$�OP���Otʓ 2��J�"C9g>�p��4>�*�k��h.�O��D8���O��$�� qbh7-�w�d�6�ĺqB�L����O��$�O0˓/gZ1�Oa< �:~��q��� �pӥ�&���O<�O����O4�F�O9�bUD��H�N�D�F��%X���I�T������I�k\@��I�Γ2T.��5��HF�s��[�1�	џ&�4�IQyҡ���	:392��(�� @H8)@�����O����<���8��OK��O�����EE!09�ij�k��tW�ȱ��'_�O��;��꼛ՋXQjPu#��R:��D�G��P�	����5�����Iԟd�	�?��I�#��m8��m�#`�qbc�L�D�����*ӘI	4c��>�!���&�-�$te�M����( '���O$�D�On�ɩ<�O
��r#��|��fL{䐃��'�b@Y�.؎�h���P�	��<�1��ܜ��(H�.�//��̰�J�I��A����	l���Z�iˊ�2�y��ߟh�I�XЂ��}ob@%eU2)�d4v�Q���A�I����?����C&2t"9�����ѕ'��'�ayb�G���9 Di��E$�3�[;~�6mX���͟���^�IƟp�H͂\Gh5a c�4�"����p�fie�Q�<��l��IQ 'hH�bW�LX�t���J��M0�+��SvX���A
!��x��(4�ZXZ�@k�pT�#h��C����Be�HPc鏡u�!����q��سEKQ?�1�@��k��ŀ2��6M�L�P2�����kZ>��8s�H֍+�D����K"t�+�A���Y(���Z�[s��t ��'����?����y�	�?�����tG%�, AD��n�嫦c��%���ʹa�Ȕ�[�N_��-1�/N���<�h�1��(so�0C%�#�+��.^�)�n�1M��/	2R7�8YF
�O��{�Rm���G�Rͨ��K	�E2Ȝ"e�IhX���á�V2<�dGՙ2:>@�"�%D�(Q�\"
kf���T;h\Hz�!��j��IIyrIB��\��?Yʟ�xx�	ٍ0�G�E	}��-͝��'B G�dxa��2A�m��g�O�S⺋�$LN#��u��ac��#3��X�� hZ� ���	�D�W*��O�Z��i��*��W`��?� �`�}R����?����H������'ʺ1£��}�Ha�.@H<�#�0"̸BV�X�i�:L��AM��(ˉ{
� ���V��-ax<Xf��*q�L�i�B�0%�P��4�?)��?��[�xx���d�	�b�c��G�V�cRIR� 	ԁ	�NN�2R:		WoѮ���^��1�>��ĈB+DH��؋��� #^b"R0 E�X	r�P9�'�"}�'���T$݊a���QF�P�u �� ��O��+?���~b�}�)ރs����(3��VY�ȓ-�άȷ O)j$KB���P\�=Y��i>������BEIP�f{���%'��M<H1�⚭�?�!��s�Ȼ��?A���?�%��L�D�O7��C�@̹!��M�f`z#����M{��_Y�Dh����|����2gb�����x�r2G���[~LnZ8j����ڗP�"��"�V8��3	'r���.(|�Hq�e��-�D�'0�X�I�-$*u�&A��yt�b�A� �0B�I�6�����?`�2��4Jr�l�<��T���'{�q������ң�UeDnl�gӞ&˔�#3@(�?���yrBƹ�?�����d��H��PFE�t�Y�tOP��8!r��L+	�lݻԲi� ��Dۂl{0a��o��m����p"J�&,���(ɾdk�rn��	Il���	�dL"�'{���Ֆ촹zď�D�j�:%ǋ�(O|����~n��I��z�����4x�!��S0�h'E�%r������8�.�ʪO�=�b�ꊾC~��a��عkL�taD�VE�<�%��A~n$�p�Q�xڔ����i�'�����FqpЀF�5Ĩ�*Oh	QSɿuv�!�w狕U=dp�t"O� �!�ۮx&T���iR	)N��s"OR4:�m��P� ��Ի1	��A�"O~�è3U�\:6��(g��p�"OPف�B��$���'�"�ؽp�"O�%(�.�nF=8�A�c���"O���Qi�	I�V���\�r�F��3"Ob�pB�7*�Z��Ům9&  "O�qT��	f`��OˀoN��e"O����*A+#p��Dh��Р��"OP��u�� ��QW��dɾ�1�"O���7�˜z��0�EFԤP�a�V"O�ࡖ-�y$�a�%���##"O �aЋQ
?����Y=@�0��"O�I�*ǳ8�N���O�%MH��"O@1���Z1��2�G�)�X��"O�	�w�Y�:�0DIR\�p"O�(赣 #{ �����Թb�"O ��'��%Yda��,J�'����"O�,ፄ�z�ѢN�up��F"Op�Z�FV���s�֙<v|�2"O�p+�>3�	��^;����d"O��yEFX�pE�PH��1��Dl<D�d���=��D!�(W���{�l=D�|�� �-�R�+%�D�K�$Rwc/D����O��wa��b�dB[S��{��/D��
���9	P��:��&h�����)D���7 ��u�>eR����t��"D������. �,\��J�`��9�� D��	�Kn�u%��<2���i!D����Eٻ	=�z�6ʡ{v�!D���t$, J����TNh�XU�*D�LG�5XtN����}�Nؒ�+(D�`P�Ȃ1y�0�CF�r.�{��:D�X����8w%y�̙��2�zPL8D�����>DG�$�4� ��!�#D�h�� P�O���7f������ ��`�� 0�'I����m��q��
��$͇ȓ,�B���Ьg Zԃ�	�5�@)Ò��:*�rN>E��'���1��B�H��I�nH�<
M�������%��4�� ���|�INZ�r�M	S�a{��
 J����b��X_����T���=����"X�K��j�6§��\��a�97+�DD�<�3���yƬ"B�	�w�&��х�C�3��P�U^8�"}� ( ���� J8�A4@ŚO#f��S"Of�ڗ�O�t>tx�����G��ԙ��F�x����W�;�g?Q���r�.�"���Ԥb6kq�<)���<�H��D+ƫ��@�`Aٟ��7��	M�v����'��[��D�n/dh�t�F����Z�M�f\��k�*6�7��  R8]U��)#��ʠ�V
	l!�ĜVQ���7b�Z�vU�O�(�c.�:��$B���H bvNX�0�%o�����I!���8|�H5��dڜSC.̻�fߤ�����mI�ťO��}�����������Q�Z�5V8�ȓ)B�R3��"R�L]�3
�>�m�I.4֐0��>�a{��Z���-P�+52�f����}�a|�)VJԵ��'�8����]�a,N�mt��'�б�����U��ⓗq`bK��ְ�Թ���ɗ�w����-E2���je�P!�����Cv)B��mib� !�:-�څ�%�]�!�����n�<2�!�$Ƴf;[�%���R�p���.v!�d[Xꔀ
EOX�>t>5��8�!�D��S�����bV+8� �,�># $+��*���?!>�)m�4S A�9�y��A]�K� l��f�6]��m]-g�(:���J^��"���Rf�!�OrdB$a�)y5�D��0�Z��t�'�n ���S�=g&� #�Op�곀:��l�a��
va�9W"O�1�2F�*�Ґ0���u���t�xB��$,-�D���;d\Q?�as�S ��qG�A���
U�2D���%ڕf��b/Z}�r��n-T�AAFQ�����J�����q������B.A�"`�p(Z7[L l�ēt6�A�C��]�̲kX3:����6:?L���i�-�p>Ѵl6}�]�'�R/p�t�"c�[X���4K�X�ع��FB?V$ǋJ��e�$F�	�،Q5��j�<�w�ͱ?��(�(�:�H��_��<|W�]�1JS�;�F�E�dIY��`�@�L��f�||hQl�'�y2�MG^\#�@Қ!���F��&Dn-�$��uyR�2%�b?OVUP&K^�b ؜*PEG!0+r0�Ofe3*=O�&��bI�
z�py�B60�8����B����K�>��)���Q��� h�B]�̊Rn�-0az"B͡/EbM9�S���F�GҨ��fQ����Il����	k������i���"d��3(}��5Ɍ<_ayR�B�dW���+�Yy�5F4�	7�׬|1��t!�y��F2R��yò$@�8{�\�3��ēu����'�?������E�PP�F�ɛhֲ��g�Ia�<�CJǞ%�bx�G�\�@�� :�iB=�~�Y�	�{�̭n��F�*}�c��<Iў��g�܌?��pDJ�sCШ���><O��P�P�qAڴ��Oޟ|$�m��`�!qi�sS��t+zI�E% �.)B�&Nxx�T*F�/HE܉��䙕:Y�	y��;��I�)s��+�j�O.����Ⱥ~����K?���Δ0�p@kޱ
@������ !��Y#n��Ԁ�H�#;�HK��I�Ҷ錎M�,�)򃈶0��p��9��Lx(`��wV�-�4��)%M1P�ٸ�U�'Вmj'�İS���:.�v�6�����v�X4S��K�V�F�p7M�F�S�,ų�hOZU)/V�5�Ȉ� �#��`E�'���`G��T�0��ƪh����R�( fc��`	|`�A�'�^	�+1a7a~R,_#�~��B���kd�˃���	�%�H�ŀ�K��r�Tx� _���{=��A�C�TpQ-
B&B�	�"@��hB�59��EY'aE���k���
$P�Q��v��0�=�)�t��4�}�,�u	��L�d�d�9Eif40bI;�O�!�%�?n������C|��� �Ht��'���z�@�y�����>{g�-G{���.S��˃��/��|��,���Olx��.�P��P�䤚�b���Xd�7�-[EQ8ykFT+GZ}���A��Z�P<���k���JF/���� xG�1�'�hI�s��[��طtzB5�)AC�`�!�'�|�&Z�o(z��v
�3����H��y��$v�l�Х�������"�#C��x:gɇ�_^��ѩ�(`r��~$Cӑ?7H��8�.�S6��6�k��Tz_�+��'�2�{Ţ�<!�gB�f"��c�#?�I�aE� )��`�炽t7<����62^��� p6�s'�#�S�? ���'.�2<�f��!A�*;�	�ƗxICdP|L`�'�z�GR'�* �F7���Ϝ<!��ZQk�{�v��GL����S��ͯ����I�@l�M!3d�@9 Q�0!!ۈm �~ӄ �S��N4�r��Z2
��лrFH�?�|\�ā��E�ϻ u�|��DvU)
�NR.�d�;E2�2��GH��x��tgH�9Յ��c�|�T�юVy�AG�TUU\�bV�FK��E{؅��Օ�y�(�*cP���u�(ųD̒�p<��.�p�I�D��O$0j�
Xs���`4C�+ɾI��Hݏ��0`�N�C:����l[4�M�B�У>��(J*t��D(!r�p{��W�d�SH��V ��?	e)��a���H�DO�m	i��%z�9#�?�zS��U<ThF!� +D��3�:gM��k�$S�5�h����]�`T(�I?gO:QxÈF�NwʹV�Bz��F�q��ϻ�b1�G�/&N�e1�Ō�Y��Ʌ�C��	@�D� J Аk��_�.	��̃CAj8�tM�����A�1m��(D�I$Ԑ�?Y��	q�,�����
�U��$_o8�L��k's<@F�O�"a!�s������"C���r���G�w��(IT(:�}����+1������&�%��3�I�/3"H�'�(Lxw쎒7XjH�OP�����%%Ҙ�h���6 �� �'���gk�-z��Y��i�!�	��-!�DO�!�
���$! U�Dy��p���D.`���ڦd�iA!��C4���6.�j��p�݁3!�D�4*oؑJ��R�y@8��Zu!򄃏.�}�rmχJF����;.!�$N�sU���S�5[Z h�
J.dk!�l�$�5���h��)W	H!���6e�<�x�N�:j�l�ň"�!�4��I �?[F�8��N1=�!򄔯m��`S&ċ�v�!��-�!�$E�K��˴��,Ӡu
���	x�!�dH�A��ѐ��-B����B�m���~�	�YG�eZK�(sP�z��^�&~\��&>��A���<��6$�B�K�L�!�6P9�ȆU�<��?'�`�p-�6b��a1��S�xZƤ��$O�~���}�BH&��̪�f."h>��OJx��
E���<	��[8l���"̒�H;��8�+ɂª��� �.��ɒ�H��ɓ�̹&oѯL�n�`MW���#=�U	S�X�}*s
��C���&Τmd���DQ��i��ܲ��ر��'�h�:%h�h����F >Q�nݴZ�!�b�2�)jCm�z���(FJ�O��;7�]�&*��أE!H�k7"O�D� h�&3٠��GK�jM8P�uU�����Yf�XC���-j�T(�'ZTЋEKu�	�:n��!Ð������R�a}�-�;$�����9ia�������YCM/@"��Ӷ� /D�n�8o�}�EHDy�O ��+�H9�b�EI��q�AX/R��#=ٔ.UG���}�0��Db0��e��#�q$g�� )aD�C���̙��<�êf�B��I+�a�q�ă���b�
^P~��dئ�H��'!���ǃ��MSW��~PNx@ U0oE���f�Q�	������V���
[��}��G�?X"D�@۬Ls�l��)5��O�z�\�h�� v�d��W��ب$NM�(���K���y��3C�`y!TnB�#C����ݻ�ēB� ���9t���� K$RT@'#DN3F��Nb�<y@��,i��$���VW�D=�IޛNF؂N��R�G�����ē81�ϯju����/��]Lt4�ēDE�t�@AY?b�����a���T-�#�I�	��f.>�Oi�w�8�&���ʄ�b��'p�Yz'aÕ
 ���'\iY�&�p_��A�̓n��Ļ�'��X	6�ɊKGf�A1��c>��L>I(Za;���'.�� �g^(���9F\�5 ԅ�(G&�8�$ �x��5 U��}:T�RD2�Ɏ?."|�'�f�CK�����r��7�Bh��'�ƙ8&��0�`I��U$��I��'٨��!�@F��qXю�-a&!:�'�y�SLγC�0@����XP����'Ж��C���Δ��#�Y��y�`Ի/�����EN4p(4C獑�y���*x<����4��A%���y"�ߴ.6�tKq����hp�C��y
�  ����
 �P,Z���H�"O��@޸a��� ��ڽ_��Eia"O(�Hġ�,'�"Su���G�$S�"O��:s�+��PeM-
9| �"O�!�cJ-�j H��E1C$䩫�"O��1cL�f���hW������"O��!2��joG.���Y 	�1qZ!�77��8+6l@4̅8F��42!��R�d=�#��B/@�v��AD"O�؁�l�14�����L݊X��\B"Op���޿pԠ1x`*��1�@"O<�K��Q�m��0 ����4�D"ON]���ʼb/:���"�Pɂ"O�I��!�.]���k�H�4X����"O8�h��ǀ2b��Hq�	9G7�#"O�Db���="H�p7DT�|8�p"O�9r G��FI�U�Df2 �"O�Q����D�$�/�8R@"O��3C�8?�1�ЫK�g�@�v"O(��K���i3d(X��92"O�`���^o��Q�ٙz����"O�l"7��4xЪ��Ŋ)s$	�c"Of]��n�GGm��H':����#"O����撵�7b���쩩�J�C�'�J X�/_Lِ��ËU���)Ox�7��'�N	q�/GZ��T9"O6�y1�Λ40��:�#��@��"Of4���Z�0�h��7E�%q�"O%�Q,��J��sǅ�	rbyX�"O�8�C��i���f��6S����"O��CU���"B���ŃGnZ���"O���? *�`���1�t���"O��i���\2��rEW�D�J��2"O=�'B�� 8 ���BJ8O��|�"O�sE�D��AD��zhv%	�"O(	� �6)y&�Y�oϯ���#$"OD!�C�A�L����IR��r"ON�C���j�r��GÅ+�@���"OTr��ܫ5�"���-D>��چ"O��x1�� �%'�
g�H|�s�H��y��
�xaL��Z�e8&(Ӣ���yb$[�y���ZR�0m�tqP�c��y�BJ$k�z�ʍ�m��=3"�$�yR��2$�~���%iϸ$rbj��y�a�8�$���c��R�Y9��y��/X�L�*�/ދR���������y�kܦN;� ���Л�|(�A�L8�yh�.�\M03K���Y��L!�y�e�w��d#����&�.�ybiɄZq,I �g��(Az0��)�yRgI�2��Œ��t�P|�j��y��07 `%xq�ĜhY��͜�y��IL�X���X!b���QB�4�y�L����Ձ4��[�n��BӋ�y��S���`�+T���v���yro�pt�9�3���B_k�Iչ�y��W�#��a9���n�(��ٽ�y�˕�b��J#���9:�H�����y"�� dp$y�h��^ ����%O�y��
 $�U�I�.UHV��)�/�yr��;I�=p��@Nw�U�Ǜ0�yB"X�]zB��P*ʗ[MI�D\�yH�4l����@H=4��vX��y���^P��r2��(��(K�䝩�y�f�a`��A��
i���ZEݯ�y
� ���TO�\#0mCԋЫl�(mY�"Ox�Fd] cĎ�6A��6�����"O~1��8A!��*2C�zh�X��"OX5�4B]�fI�)+5d��3R�����	�"�V"~j�� ~������^�
E���I�<��b�v/"3�[12�9	��<!w"�s�����HB�	?yp��fI1�
zP"O�bG��z˴|���&TՔ��F��H�2�0�O�(�Fb[2�a�Խ&�![�'��A�'d��	��D�l �(�j�^$Q	�'���H�k�ꭋ��		Qx ���C�?�?�w�؏.�B�ۡ���e�̐���>D�|����LtD���G�tj�c}�Ȁ��!�S�O�N���k�<&�@i�⭉5�VHk�'���0�,7�u�a1Mp��O~�B�'��$�w�ĠP#�^�&:0|�����f�fh���Ȏ6&P��H4����{[	BgDX��x�@g٘*��G|�o�!ň�ja���'6�(\"��M~Bk�"Onu�&��+YǊu��ڀFf�հp0Oژ���)�'6���c�ܒy~Ҁ�r?	�҅��wHd�
]/Z
��]<tQb��Oa��'�&��6��
4��La�� ��X�'G�!�%,
�K���ff���E��'�^���E�a'�D��&I1�P��'���JY�8Y�t'�����'v:���@\4f�$ s!I����в�'����D���:%��Mܟ
->\1�'��p���V�Bt\".uVH�'r i��G� ��0�0�\(�
�'�f���)ƿ:Q��1�5���B�	!mj��5�1yAh��b�F�:��B��!LR��I�G-iL,�Y��^�ת7M�:=�������g$��2�%H�q,x���ٺj���$�+���'�y�ED�]�j���DMLK�|�'?�!e��7k�T�g�˳@g�L�}r,�$��i��,˒@�����8�jp�A�¦S!�
#*ʼٴ��9�
i9pԬ	�0q"�dCz����×6B��)�Z�9�J�xb�N�!��;�pL�Ԁ�޽����R�!���)�
��l�81y�D�(:M!�L�>d�;#���<xD��BIQ�A�!�D��N���c�ٍSa*�K�%̟n{�''�UFy��h��T8�� ,b��rA=�y�Wt!��+	"4�f�B��\P0�@�M�@ �(R(�.䚍���|R�I:>�r���F�z4���b׎ΰ?�ա��4��p�2D��3�� (0m�[�% �h����w�� h�m�S���$ѠL��4��f�9.�n�c3cٚ���d���/w��p;r��]��LHhQ�n��'&H ;�<e䞤��5��O�Ż%�Q}'��S����U:�3O�s
�����gcF�g������Py/��?-�Q�ےv�$�@(� ᇏK�!��ȋ} b�s��<-�4�.Z�W����.��5/��ƇQi"�{��?Q���a�ɺ*F����*� P���G�`[���W� ����f�Q�Oi�XC���>I�8$ƥ!`���
�``���d��GJp|��I5W�Z�� ���[i�1M 7��=iVŅ�V�0��a�N�LaP��ޏ"�Li*�R�Zm��Y��AJ�pe華���ֽ3N9�&@='c�X�����v.�	����h�)K�~�y���o�2��LB���c��Ai�Y��E�\k�l����]�<�B�L7�~���F� �c�.O�Z�3c얞Gn�"2X ^���O��x�KS�ɹ��A�9M�0�05��_.���d�?\;��D
A��rUH�+�J�q7A��0�����7MdA���s�Ks�'}��@FO!Iİp�Iݨw8�����ԝ~v�H"���D�ع�"b�	x@����É�i�0�y�i!b��0���:�jT�B#���`,���azQĖ�jL��H�&`ӌ�x������Q��yaN%���A�s��(��S�s�� ����)X�I�jI<^_d���"O�X2��BNQ�=�ABӣ;��cTL�3����ғ������)ڕG�Hixp��Byb�1Q����܈w� �����>���>�.q�F��~]z5�Ly�M�m�+�MK.Ο+of��'��)²lx��	m�'�$AI!#�=#���Ӏ��
�j���$�h�de�cl�ڰ�aRMNaRH���1f92�S��/��Z��Y��p?�fܞrZ�x�1)�if,C���<)�-�Z���b��t��=�jĮ��s��K0p�)N8>����A��->�l��XO&�"�Fǥ^�����݇x&����h
"��]�sZ��1`-�t�X{~�|�g.���r�!�?iB�Ë.$ Q�2�.LO$��aEP�I18�"��L�	l�;a���K)�A,�.�@�Z�̞�s�����JP1XDQ��	��G,4d�����6~��iI��,��4z��I	2�|���dhJ��te$�Cڣ�Ȭz��Q�Ѷl)� ��>��<��'�y��EF3V4$�����Oz�Yb��Eܓ#�Nr����O�B���)�G?�qfhޑ���S�Nl�i���|:b�KBM&D��8���6�B���N�U0��5�_�'�HHP6&T�\~�YT��<�BN�����?ARNև$����5o�m ��z���{����F����.��ѯњWH��ÏhG��I�>MV�A�7M�~E96�'�6|��fۓF��c���/��1��66>�qÄ�M�~Y82'҉k�48B����v� �����c�"B�	c�^h�Fj
-����RCʃ9���<�c
<#^i�Bb*m}�c>-ã)@�a(�xS=�|�0s�2D��їkB�jM� E,9���s F?=91"��ƄIbPŐ�Z�z�`"~ΓJ��Į��:�]�S�ٻ"�t �ȓZvx�kRH^�pu��'K$�"���f�D
S��>12��C& ҁZ�x�E|� /��(�"үK2��檛0�p=��#Ҳ}���"Ă3\��yx�GX�Y�r�AV��]��1� ��'�����"�`�ܡ��hTHڵ(�9���C�����5�=Y�hJ(S@�F�����;0Lڟ���� �u��8���1�#�#p�����y�N�&�v�@ԆC���Hg�\�P�uiFc,�8u�5ϡ4��_�b<f��?�i:��bǏkjd��!�2�F��e"Oصc���%8���ȝ�W�.�%�m�x�#o��<y��B0rصa���xz����l�	K�H��f+��k��p�����p=��%�\(2Ez�O'0H!���B�LU��� hH2$ʴ�{i,E�P�PO6�-,S���<y�,���ԫ���$��$�^`ܓ� J'��&t)��N%7>�$'�$3N�j\*h�倗^���lR��x��W�Pz
5	#�CI/�	Y�a
.}�x�
��@�pr<��𪋰e����'z�n�W��D�jÿov����� K=!��%M���rp@ؾQ�@�H����M0Y�>�$�S�� �G���A��d9�I+*H�!�t�I��ǎV���DJ�5�v��$�,U�z�ZR!��zR�}ZФޡ&
	J7��e����#�ɇE��h樀�4�ax2倊SD-�d��.R	PT���HO���vH�	be�TB�D�)�Q�l0�Y�E�P��e���`�J��Rn�&sP�B�I�)����E Y�R뮡jA�T&�6˓$�J�������)�h��'�~�Ş@�T03�"L!Q�rB@�-�T��Y]�r�;7(a���Xg��э��og^�q�
�<�q���|��S~�NW$�I�$�~�٤*U1�Px����j��&*O�;{:%ڣC�5�� HĤF�("򕹷�C�}
0�Yw�9O e0��D�,X��b�./N^
�'��͐/ޜ�(�L&���hJ ���*bޔ4���ӳ��
ސx���ʔĳ4g��w��c�m˿[Q�M� \��	���/����Vg&%��X�7���wp�u��,�&h�"A�'�\�i���
�'X6��G�+
��s&ޞ*
,u@�m�
��4�'���B'��G�)�3?	c_�[�F9𧅎(��$A,@���5&Py�KЭu�ƅc�:7��QZB�%mڍ5Ƅc�F�����	�<�4�!�k׈p��(KPF[Y^"<i�#�	��%���O&���
53]�Q�R&��u���	�'J@I!��O�Hd��9)r	&��:�O?牓2��d �Y����@)��T�hC�I4B.���Cѥ��8R*],C�I� �li��� yX�9�1 ��O�C���(�ps�C�LnA�!Z�C�?y���k�<5Q��@�w���K6"Ov�A��"�$C	�&A �Ƀ"O� �M5��(��P4Hk�v�{6"O���*J�Ra���f�N嶼�V"OX�(��+`8��Q'�ϖ-��!c"O�����M0̜bc���:n��"O� ��2;]�4����i�\��"O�őP���v��$��E�;��;W"O�T�A/\*��1�qeO0+R�@p�"O��+� ���nߥ^O� 7"Oj����L2b;���dސk3&s�"OT�R�ōs!�w#*0�,�@"O�*�Ӏ?^�5`5�� b��"O����w`Dih�*Q|2:dA�"O���V�:mC��J��<"d�"O4��6�yl���$�2R��P��"OB����x���e��C�p)Z5"O�p������M���ܤX=`�SQ"O��k���8#Mr��ckO�0;��"O�U(�b�~$���d5��!q"O
x#��0���午kP&�Q�"O.鳲mQ�4����PJ�Aڗ"O�"��Փ	�<"$LF64�P8�"O��ك�[G�4ĚPe�2_�TYc7"Op���9`�=�Eb�=y�=x�"Or��-��T_`x÷��;)�h v"O��Z�-� ~�2��@O.;epU� "O@���#�=?�6�*'2����"O -{�5*m��G�z��u�"O��R��N�h�b'�5� ��"O&"%B��h�
��!�/+����"O�]�@�BJ$��1�%�C��M	�"O�x�o�D����R�T��h�`Q"O�D`Ð���sCڃQ����"O�\م�M3Sr,h�뎮Jr�@�"Ov�#g.6-<͛�+rԂ"O��H�k�ton��C��0Z�h��"O�`@d��y�kƿ1|��rg��\�<�fbwǢ�
w��&cj�}���EX�<A@�$M~>�y�jN�i%� �ң�i�<)CH	�t��ЭJ���� b�<�4L O�L����C�jq����c�<���D(�c��X�,����B\�<��N�&D7F�а��PͰp/�m�<�@��\�>�n�5����H���y2�f�r��R�O�-���F��yV!f ����u%h:t���y�3FZ��0G��fHVLCӆF0�yB,��{9�H�"��8d.z�aw&��y��E�zP������\ܺ��K��yb/	rdJ��ן}�n8��*�6�y��36��x�v)�8sZ%KbD�(�y�M��X;P���k���bƋ'�yr'#"�.e �)ȫc����N"�y⣆*�Z��G�\+�bS"��y��,ibDƠ8&�a(2ʚ=�yr?��Ѱ��*���b�y�̑r�@A�
�&�x2Q�4�y2J�hĦX)��?������y�BT��;�?	����P	 ��y�Q-=R�8�!Φ4	: �ǧ��y�Q$o���j�`�'��JrL���yb���>����b�A��`R'�9�y%��'��k�/n�fI��ղ�y��A	b��T����icJ��ǉљ�y��
�%A�٫]�ҙ�1G�y
� ��I�]Y��&@^�*�t��"O��1a$;�j"�	G`#��� "OJ��B�:�x�;C�^T��k�"O�AkWl[�f��P@�b�O���C"O�P�F�!74�`v��N�fԫv"O�=�% ��hc���J�j��թ�"O0���-��!�t�WJ߇�>��'"OLiI���O�16g�� �X8��"Of�P�J��>����,�g?&�p "OP��d�4c.�X�J]3�]�"O�%(��V�;���8T��8-tPK�"O�l��o@!Vi*�t�ۋK��1!"O
ALqIh���	^��GGա�y�)��w'P�@��X���� ��y�(�>)�K#��L:F��bɝ�y��H�ԲT*D!Go�F��y���	���	a��FSzM@F/���yb�M1�6u(� �EC��5�y�����,Is�ءP��M�pM��y����'~�*0�O q�=�����y�-\�j�:�t�ʻJ���0��ybL#ڢP��m�;8��rp�� �y�͔�Q��݁A�X
00����y�!�N�ԑ�AY��%���ư�ybς#'�n�`$�&�$a�FFK��y򡉲8��ݛ�AG0*�����6�y��!lD�}ذiׁY�X0�c���y"��8�R�x!mD�#$�����yҁX�1+�d��ەs҈�`ٶ�y"�\�`����?���BH��y�Õ!�(�HH>�T �G,R<�y"����XY��̯�֕8��A��ydøی@X�NS�-+���y��G'��(��خw���C�����y2�97��|6-�"D�h�c&B��y҂�42�9�Wɟ�FE`��Ū�y�BV�8|LȻt	�����⌗4�y�-��;?č�S�ʟx^�Yud&�y��G{�+Vj�? ��y�����y��@��ԝ{$�]ۢlS��y�JG_]q1��F�FsP�����y���8u!$4ڱJ4h�씂P�0�y����b��G�I�t��G��2�y��G%,\"�K�@�I��(�y2 ]��a"B�;Ȋab�oһ�y��$UPְIJ۵6�� ��#�y��;J����	�4��ё�N��yB�ۯX1fE��'3�b/�?�y�+I�3�X�1I� ߂�+!�O��y�C�B��fᑶ���a���y2�
!��E�@�T45Cd�i�����y�A���ۓM~5�wE��T~l)�'I��P5�wrW#">��)��yr(�	�^��U��4	�3�y����R,I`gF�GV��b����yr�G8A��p�A(*��0:�i�<�y�b��8�e�Tn)w�.9GGݤ�yb�=�ĕR2D�)&7��) � .�y��H���E�&2��y���3�y*]80}:�p��;M���k�$�y Z�^��E+� ٶ�Ĭ�E���y���#u�2��@>Lo�03�˅��yR�YGf����ꑍU�t��F��yB�K�,����P��t &ƛ��y
� ���v�����+w��a"O2�iq&�����(�%���Z�"O�����49�����F�>t��'"O��� )�}�ٰ���M>�0�"Ot��q��v�����]�<x0iV"O>YS��]+�B���+N8�y��G�2��Ή�<4=bWm���y�H�aYl�֣�,l�FaT'6�y��'?�!��G4PΊI
����4S�C�'8^� ҩ�?:���֪0a�6%8�'�HтTɞ1 ��	i�CX5
�Z�'�4сQ>n[�b���4��'�R�[�̃<�����	)�5�'���
B<Z<(鱆Fӳz��у�'�}��&I�q�6��4'o��#�'�����c��gj�0L�3�'.:��/��0g�e`�.x��'>����/\a�LE�>r�l��'jf�2�k��0�24�4�̢j��s�'
t�XR�N&PXHsB�,(�X��'	��r�B�z���7�ޡ#����'���;�C��!(�S�;�`��'|�td�r���Q��  uv���'~��9�K���� K/G̱��'��]
�ɝm_�#��ıP� �';r�ї�T������Jz��4�
�'�8,ؒ�әp}1�	�x:~�a
�'���J�*'L}�C(T��.���'|d�,�$c*�9��޽J��E2	�'6$9q���Q��9HšH/ 0�B�'>`�)��X�[2���^#$�D	Y�'=5�"S72L8�E�Q0Q�j�)�'��R�FKX2E*ug��O*���'[�Ј�A>S���[WO�h�'�����i�>k�H��/�H (���'xҘjU-�D$ F�U�>��e�'�p�ȁ�_:�r���X�7�|���'��9�F�!#h�=X�j�z���r�';|0;�H3Z�8�#�Y&"�n�P�'�LEB�%�<6� �b$PQ�r���'�X��N[�:�ͣ�Lt3h���'��� �B	��+l�p]�	�'������\�,P�1���`|px �'X(,����|��yaeԷq*���'!�Pn��-���Aw}��H�'�f؃B�K�	(L�� �|(zd8�'4Fpr��'f;��a���`*ج�	�'�J�����?M`��PW�J�p�'�����
I�_AF�Sh�w�0��'߬�;�,H��i�c���S�4��'�b|��N�+?<"4$��
�Е��'�&t���ń
a�Q�cES8{��Yr	�'�j� ��E
{��)�.�!w.���'�J ��*����kZ$N��@	�'7<9�D�1�Ĩ��EO�s��	�'Q�A��A�>٘��em��q�'yB�� �3E!��J؊ ��<��'�rt��&�K"p�@�+ ��3�'�����m�	\&TY#
� d���'�b�oBQ?n�Ycʋ� ����'��u�D&,�r�iѪ�W<��'k������> ��`�0a��2�y�'�vِ�V�j=��(����<�P�'�:�����/��,Q��-F�9���� �4p�P�\� �"�Kn4
U�A"O�{�gE�LF*�`��� T�y�"Ovh IP+o�T�Y��rl�}�"O�-�#�s1� �v�D%��d�$"O�xF�҈���� �M�nέ�"O��8��<��ѱ��rb�S�"O�yQtA�h��%�����]��sb"O�С���l��%�PA�6AS ��w"O�u��ɐmb��Kb ��C�"Y�"O0 ���S�5~�Ѯ��.�~�ا"O|�b"J�h���N#N���)�"O P���S[.��b��ߓ�M��"O"h�[�����?6�y �'@��y2e,�~}1)�@^ep�A��y��g�����1F�^0č�*�y���*I���B��;O@��A�y��R�.<� ($�-�$�wgN��y�c��rPd�n	&S�a ��7�y�7D����F�3԰��R�A�y�̀6�E0rM�'|�l���f���y�cVt� 
�Ғ��INb~ͅȓ�V��%[r�䩸¤��0����xJ��/��7��,H@�5_\����^�y���: li%�ճ�
�ȓ+����2f�?0K���4�ر2�&��ȓl�`����E)��( �ʫo�8=�ȓ�aA$*LDԜA���-�q��:�p��ʂ�(�)暞`^�ȓ<]X�P H4��źV�޴LF�ȓ^~����%Y��
�	21���x|�#�����iR�)��̵��tYu;B��~6����\����5�z�#k]-9�t�CEL+&͆�g���� BY+13������?w�,��$�#��ȠZ�E�QMѻ��U�ȓ�LT����غCCŐӎ8�ȓ�P%�\,�`�:��W�(�<��6^�a2���>	z�kc��	HV=�ȓ+l��y1��; 2�EK�/�f��Յ��a*��ڱ	�L/Q��hHB� D��Sf'R�
u��j���8�Վ?D�英$M�3@B5����1�d�'D��U%�R�	�k�JO���.:D��)��+5����M��WX�۵�+D��`��������N#C����*D�p�TJ��h�p�Dڦ��E*'-D��ŋ��\ͺ�&[�zA��*D�t�bKV�n'B�Fhƴ�F�
1F,D�� ��Ś_�����~�v��&D�ܸ��&x�4T�P���i��U ��$D��*')]�p���PA�f	��p'�$D�Ȳ�Ƀ�HJ�d[�+�3}��غd�$D�����~�H59�l�2Oe�D;��%D�P��j�1=N�2։۬}����.)D�0r��Q�2�&��6��{��Xp�&D���>�. �1�������*D�x"5�;�=3&獋Md��2�6D�jڽ$�;C�I;Jp8�E5D�t"��_=�H������`�^��D/D�x�*�/�H���
�m*�Xk&�)D�$�&9�K�h���(I�%D�,(�#�]44#��C�.��� ��6D��x���E2
��f¨0/�Г�G?D���G�=G �y �L�(tH��2D�� vM���D�n��t��-N3X���"O�{�V�|���=�*hz"O>Łա�;w����ǫ��wY��""O��ce�<��y����.0�V"Ov4�s��7*��ؗ��&��c"OHe+���&-�l4� �,(��"O��d�2�2����W�L;u"Ov�`O�W�����S�$m�"Ot��CY:
���BL��m��H�"O�Y��	8
�R�	��
�-��1�E"O�yӲ�ɿ9�f�h��^��<�'"O6�J#̀�0��1o�E���"O�U0��2���L	:I����"O(�;�N0�*e� FY'),�숃"OP�C�Jcx�Iz�'��xx&)�@"O�� p�E5J�B�l_�2d���"O�YXj��fY�D�$�˦cZ���"O�,2b`�
��p��
ϕ�f�j�"OZ,ab@/����҉�#^�МA��'�'����?� �fg�+V>fH��'N���t��q�]�7��R�)�'~�H�F��1�e�WƉ�6K �'���ӊ�/ LU{�GD�\΄р�'���#�@ߕo���Ѷ��3
g"�Q�'z����Y�xzr��T�L6,#b`��'0y�Jd�l� �	�]��s^b���Z�&'RՙGf��H��zCʸp�A�c%���6I����x��\"�<9R��hNj�0�EǢ4D�M��WϘ%ѤM��&8!�/�U�vՄȓ":���NO����@kA?J�v��^NpXc$(ΘV9`��2MCy=T��c.�A2���U�*u�S�A�{�4���zL����$� &�r\PDyи��ȓ>m�m���M?����*�RŇȓ$����OP�<�p"�z�<<���amљ)Tb�x���)h���Ey��'C���֔�rݩWBԻy�P��'u�u#b���mX(l��&��kN�-��'|��9¬�
B@�FG*U����'�>a%aР#V|I8�`	H��`�'��)z5IK'��@�e��;�n��'u�,HΊ Jx�� ; ���'0ƙ�aO&,����;{M���'�y�����%�ꋐ<�z�'�9�l�Ql����ň%>\��'��4Ґ��c����@�ȳҌA�'��[�㓭>��|Y���6��
�'еXr���4�n���
Լ%�X�1
�'_���O
�4�T{4�<-�	�'�l�+�E��h`�ML���p�'�z�iu
��+�� �DA�ҵa	�'�y�1���R��'�F�+�=)�'�Lu�d��B��{�j� � �'�>5�P�U/ǖt�1�� �tD�
�'�n@��	�-l�,1f���Nl�h
�'��BBb ���Q�6F��IW�p�	�'}�%i�ĕ�|e���!F���0	�'�����*�:���� $C�gy��R�'t�)7��5k�l�3���_"�C�'��Tb�%�I>4*7JQX�,��'%n�QwΊY�R����Y�U/|�	�'��|��
�(J$v`A�Q�M����'܌Q3�FW}��ђ�ժ\��R��� �`@��(0)փ��i�"O���%4$�ȉS`C��,� ��5"OD�bj�:-'Tܫ� �-$�Y'"Oމ؁䆻Z���G D�ŀp"O��AM�|ꀄ�å��l��q*W"On�	�AÈ7V�y�2\��A��"O$eɷ �~p(@p��A�Km��""OJ�*A�̈v���֢Vk��'"O���Q���N��<��q"O"I��g�{�> ��I�C�@<�"OpYt摼oҺ�at��;�,�q�"O-�%1�hI�g�@H�	��	}�O`h�8�d�-
�6�b&�ȼg��A�'���bVM\�T|dq���w��(��',kf`��L��-`�M-t��h�	�'��I��f�5�8��Co�Z&��'<���ыe#t�X��b6��
�'��L`�H�Q�~Ԩ��*%4��
�'N�,��HL�w����V/V�4�:��'��h��S���eh̙�Ah0���y�՟e�����!OC�4��I�y���r$TQb˶I)H˔��y₏W�H ��A>1��*�M �yB ,g�p�x��=Zg��R�OY��yr�@��l�����f�S��4�!�C�D C�΍".��)��G�!��M;PzB%b�(ŷd�����GJ�!�D�	9������!��O'%�!�J�n���kb+Ұs�TT���(�!�$v%t�B�L����l+\qtM'�$��ɣbu\<Z�@یQ��Y�a��tC�	�����a׊7
�*�,O�~B�ɌF���^Y��u�Mc]~B�:5��5�g7-��ՈҦJ�t��B���&q��=$H�A��Ȱrf�B䉇n��u�����W� 5Q�"˚1NB䉂!��EЗ��CԢE�'iBC�Ɋ��a{b��7}&d ���*cBHC��1FV�@��_�6���Ï\B�	8WB8A��(&��kE��%C�	�zjhabaD�R�xp��	f�B�I.u?�iqҨЉ]���
c��6"�B�	�py�P��\�:L�˕	�%�B�I7,���ţ@�j�F�s�DQ��B�	4��ࡕ.X�xzB��>=��B䉯jD�q��fɉC��x�ō�;b^C�I�
�@�P��;\�PH��:��B�	R���f�v�H���&?,B�	4g�X�#��Z*�D�����(B�	9,�]����3X.�9��.d�C��*r�L�R#��/#d<��<~�C�I�Dt$�Re�.H�D�Ҡ��T��C�I'V��`Pq!^�n� ���5��C�ɥn��HD�.�!�d�#vC�	'�<��F*7:�ܙ9áؗ]�.C��6;��Ӏ�X/!��q	�c�%�>C䉇J�����W��BQjٗF�FC��#^�fe@­Q�`mb�X�j��<.C�I6-�*s2�I'���B	H�]E8C�I
	��(�˓0K�SD�<	4C�U�}9�8^��0��,��H�JC�N��l$	�+����Ф�)!�C�I�o���!����f�[ Y�~��B�8�b��UL�$�<�ӧRi]�B�)� �����v�1�W��2C���2"Ole�D���
�� ��!��`�P"Ov��G'Y�2��1� � .6Eg"O,��,�@�ܑ���)&n=j#"O�d#�nC^����A��	�6��!"OL��ȿk,l{���'8��@"O|��g�#E�8ʴ��=y�X�"Odpy�		�I�C"3�:�3�"O�lȄk�8T�d�T�Աz��x�A"O�m@�CB�x ݸ�D·?�8�%"O�1rCd\1�|u;�(Xp7j�"O�<�B��8#��Lz�T�c�����"O���/MgZ~��0!�B�,i~!�D��v��IQ0M�>#�x�h�J!k>!�oLB�!�& F�0��)N=}U!�Vz�͸���X���{�oJ!�G(T�V�@���Zf~��֋�M�!�D��E(@�zԮLK\,���E�/x�!�+Z(}�`��;u,T��US~!�|v� A��
�L`@��i!�dV�(�B$I����L?� ���0�!���..��a �?L
Q ��(�!�D�&�f�y#�׫\�v��w��-z!��V��D9��Y<M� 00v$9qZ!���'����צ��So��K��z2!�C�L�FLF����Kb@��)!�$T
1����e��v�Ţ3�ڥ<�!��t�|�*ŗp��:6!�,6�!�dȥC �:�+v��u�4G��	�!�d�4�y��C�(�V�J$�@j!�\����`(�I�a�%oY!���|�V�h�/�9s\�JЉ
�'U��[�,@�jn�B�Z&|#�9��'\9rh`t�����Cx�!��'�Z)�t��D;dA�A�89����'��JIԬ�0��2G�$��'/"��RMxAz"�O.'X���'$(�b�B�Q�z�A˽%�d��
�'[�-�ר$k��<��(��t�<��'}�C�'.=t-��*ׂs�h�0�'�X��FY�08�s�f����'ޔ�C�߁�8-�$�-W*���	�'̼ɚP�U�b,�H�D(�5N����	�'I*�c���&u3�Ԥ'{"���"OM�T��.M�Qط�**G��E"OМH��N2#H���bW9h5��6"O ��ZBb]YSk�z0��#�2O����l��D2QqU&7��-��S Y*e
�<7 r8P��)��$��Z~��	b�L�a�V�'�#{�R!��P1� WB�eZ�V0�*���&D� �LR�
t�0k��'MV<�q)#D���Q�˧K<�Hö"͏JEb�"�� D���삆#��M�5bֹY�,q��)D�4s��3�|	�D�՚Q�4yڴ�=D�tӨ$� �0�ݷ%,�h��.D��qu*�y��D͚	4W�1��
-D����F�x]"��D�Y��,D�hXPN�q����$F1M7D�P��h�֒w/�f���@k�
!򄇏N�2��A�RtPi@*���!�Ů ���&�(;������v�!��L݌�c�;22��jj� A�!���;>�� ��h� >�0�v�/�!�� �<� �L"��Y��B��6ĶIJp"O��Ad蒱9ҤQ��
�Ȥ�"O�8��ߝHC��c��<f��ĸ5"O��"�s
�=��N/����"O�!��7n��MQ��G+���"O�D��H�Sl ̸��L:~N���"O�@����m[�T駃K�[	�ղ5"O~L
ԣG.���	W��f���"O�dB�	T�XB����^cb�2g"O"�`���b��ȋ栃	��9 �"O:���ʗ�@0�c	Ōf����"O*�"�x�J-�7b� S����"O:d�c��?H)� ��
�5w�\=ȱ"O��Z# �~���3�$I��"OvD��7P����@�.,a|q��"O�층ɒ�}�Pt���ʚYAH��"O�MDgU2RLT !OmQFlaF"O\���NA����p�O��(+jLHc"O|��f���Vl�ƌ,F�E"O�a��	,`�V��u���n��A�"O�a;���~i�����(�{�"O�+0CD/f��3$ܱ5�6��r"O̰�Ƕ2F�+��'�=�̖R�<��%�U),4�3_�,N���*v�<!�:<��) A
p�.�ڗE�q�<P��6$� k�!v��i��'�m�<�F�,�e��b�|px� l�<�!%��qwH��2@�u�<� E�i�<A�Ɋ�{|r|ҁ����E�� Z�<_�=iTe�G�v�ّKͫ~w�B�:0�h��O�<D�q�@���TC�6�x(��ãi�D	"�(��C�IH�n�e`'���EƔ�C�I�w���L��l���0dP�;V�B�I! �b��+�gx�24�6B�I��ء(P�J�8��8��IZ�*B��20�􋁆�z��0`f�\t&B䉭c�^$Pri
�f8[q�3{PRC��W5�]��L�Z�dd��l�\��B�	-{�.���9bJ�	��&o�B�I�
����t�0`QK%&��B�	7a�l�ұ�["����:a�"B�:T9�#�'7�Ȁғ�]-�B��"��т˷ynzL�G`
��B�ɫ1>pp툖+2��b���ݺB�	n����Ӌ �#�,��-ǎR��B�I/R�<c���/Dذ�q�.���tB��W��R��[-&����e:@NB䉰b K����^�RĈ�`��@��B�	�Z[.ʠK+'q*���MG�XhB�	2<��s�@���� �(B�;
rl��#A��0�.AK�Cj&B�ɮ|�r�Sg�BTX`֡�I�FB�	!7������T86J� ��31bC�	'���.�:�@��V�C䉳{�z��fL�hJ��swLϙ.
C�	=S��L�bƈ�JkxYLP&x<�B�	��`��n�Ziҹ�FnO�Oo�C�Z?�x�L�6\ $�'�B$;u�C�*y�L ���$0��&�_�g C�	���iy%]�r��&E�>nF�B�I1}��h�&��&K����`���B�If�Yjr�_�^�692sę�KQpB�	�WX��I�ş ��� ��B4|C�)� l�"s��OV�j�	�
 �(L0�"O���G(c(8�bȆ�MMl��"O��0Dӡw���S��I����"O�{��ٶys��9�cܥ6��2U"O�XS&H�hK-�q#Ջd��哤"O��K1��y��K��
|L��"O(h:R��56�왻gB�x�Ł"O�C�(�� ����A*|�i�@"O4�Qa���w����� M�n�j"Ou�q%�,(�"��F���"��"O��S�DٿGp�h�A��<pU"OB9"�1M����At���a"O��3GO�I��t��G7�P�YQ"O��"��k*��8dNR�|��*V"Ol�gh�Jܢ]G�|�<�V�<D��aeǜ'o��`���.0Dp�[aK9D��K0�F+B \,���"%��h��:D�T�k �UX�ĳ�,��&b�!�<D�D��X P�PQ��&�)[��*F�4D���Ĉ�Js�M�s-1P��c@3D�Ȫ�����V|*�d�(�rHXg�3D�@ ��C�&GN S�S%{�<�SFJ0D�̉�M6v !P�ۺki:���b.D���4ʅ;�z9��� .�4ȁF�-D�`�ĭ�+h�ӥ̼Zȼ��,D����(�&<Jg�K6��*D�,��ę��f	�3a
�3 z��vE+D�H �h�.K�>���H�%�

!g%D��sQ������oH�	e�X��"D�;S�ݰ	ڙ[!d��m)�PۥM?D�0�0A�(bڠ-���'i�T���;D�xY�
��Pg � �r����6D��S6(���)R� W�.��6D��"6�χ]�6�ÂU�-��d4D��Cg�F��&BC'�|UI"�-D�RwCҙD;�5���<p�~iAG�+D�{#阏 ��2�/K/V^NMۗ�*D���)
x����
�5��9U�4D����>%@�%���19 �I1D�laD`΄ �ii1)*-s�(�D�0D���I�!n������(�m�� $D�|�欚�4�8� �Rb
�$��i"D�\�Ո��0�QѤ�.c<r��#�4D��%"��k<��%��^D�gN&O��=���#9T]���m�i(�]L�<q�K�Eiu�'
y� P�eJL�<Q��%�h��oږK�D����L�<�V�"R��i�FT̞�S�N�<��ONôԲ�%܊,���Ť�F�<q��=�~0´���S�~E���B�<Qe��i�$-H�ƈ/)0� RB
��<�"�[k��AjУd�9��!W�<ٳ�߅TO,Ykp�#�>��W�q�<I�L�P	�=�&K].��x+��X�<���Ǐq-� �t�ӮH,Tsb͓X�<�@&u�\���
�WJ�%��<�4$�o�ꘘgNF�x4k��`�<aUo~|�A��OsrD�POZ����?I��D�R���R&] ~[ �R�CQ�<Y�E�mLMr"mF4{�=J L�<�vn�
P�y��2';�҂�B�<A"���E�|ݐ�'�5RL�{�<���յZ�ܨv�D�h�܂d�x�<���K�<�ht�C�iв��%�w��&�� �|	0��
�ȩ8��(���G�'�ў�˷H݈T�|�R˴^)��(D��{!
��2N�Y� ��2^�Xbâ)D������xؼhePf��KF-'D�����>x �xjw�A�w��<;�)D��#��0_z�E�5j>l��1D� ��&�V��U���	G�*08�k/D�����hd���B��]��sqa3ⓘ�"�S����Z�㒙9�d@1H	y�C�#}|"s ���q�H� u��M��B�	Z�`��D�G�_>$�t�D,](�B䉄���FGS�pf:0tJC�7	�C��E	�BT%�
Y{�y��݊ٮC��1 ��0���0�� ��*x��B�I0}�����O�W��|��9~�B�%iU�ç@h�,U�$A����B�I�ÂX� FC����N�=+�VB�	p���ÇN�Z��p� �K1B�\C��<�ru��bf� d�^;Ji&C�	5���eF�X�Aw�2z��B䉗q��6B��0�H���@�>�B�2(���2'�9~�0���h((��� ړ^s��9 I�`�|� �$t>�͓��?	$ď��d�Z�O � ��M�)s�<)᫓�d#��q���&��]���q�<��*�^���"���bB6�a�Hn�<I%(R����'RӮH�4�Vm����'1�(A�L6G�%��]�"�m��OT�=E�ԅvD��2?,b�g�#�yE� d��2T�W�0�L0�a�B��ybܚ-�L�c���sY�i��K��y҉	<)a�����8 ��mRpM.��$,�O|�D�D�X�HS��(y� �'"O4�H�B�=��%�WN���[t�'��I�B��xp�u�L�&�@s��C�ɂC���#a��֍"	�o�c�lG{��Dh�70�v09aAg$�QY5��t��'+
��%�y���� ʂP1�5X�'Є�����>��	`�DH��q�'�ЄJa�'W�f������Q�'�8찒ʔ<hzr=�G슌���k�'[������#��#֡��.�� �'���B�ƅ1L� �"6�O�N0�', �96�?ʀ�E}���'>q�wHV�X�H"�>�61J�'���%��Rw����`7`@B�	S�bՃ���U4IA�L'}��C�a�|���"�>�A7ʥ�j���<�Ď��M�,���&4)�m�3hJ�<�7Jy� �	W��)>�R�G�D�<	���L]��+�b%f�r(��o\W�<!�ǉ�W���Xw�� �$�FMN�hO?�ɶ��M��W�y>��)�SqcNC�ɜ
��[/��t���R">hC�	�����V�� ���$%�B�I��D���$A.D+��F�h���G*5D�@Q�޳(rPd���/<v4��&e/D��� �է��(�%R�n|�Q�m D�������p����N�l�䠗�h�F{��Ʉ�o��9�d� q8Q�EY'�!�$J�4��&�U�z�|<a���6W�!�V 8@�h��3��\����>J�a~�T��zp�Z�"Z����Ee�}b5D��B���C�i��%u0x���8D�� r ��ŭNJ]3���%#nh��"O��lجt���?]�0yz"O`��o�jS�����x���f"O!�fb	� ��\YF!�\����"O��w�N#J.��Ti�"O�{��)%�j�"!��!���w"O�� V��G{����W�y��X"O��Ƀ�]�FX��.^ ]�z�"OlЫqȏ�젥�%�
?�|��7O�=E��.�
j�Q邧�  ��Q�E��y҆I�^�1�N��.�i�C�y"�N:#��F��3�N8sC*��0>H>�����K����]day2O�c��Z�v7��=�<�[5G;OТ=!%�˫C�q�U�ޯSD��[f�r�<�*ڇ	v6!�ҫnK&�˲ �y~�'���G��"V2X�s,��@��P��'Xp�b�/3�Vu��Y�<��)�'��r���Lޢ)7��%H�2���'�d��1H�C����V픨Q~�S
�'�<Q��B/r��h6C�ZF����b��y�K� ~jeaԁX�X���+�eŧ�y�M�XU3A���X�,��E���yRBj�q3���n���n��y���_	���W攞`�>������y�!-m����.X1.�"��<�y�E$��
�K�9Q��]��)��y��J��݈��&3~��s��)Y��O��3?q4I�
\��:�+�����k�C�r�<�5�E"~m�\�0GD$�\��$��n�<AQ뚙D��RqD["j���ڥ!@n�<!�*�w��*t �2okށ�ug�q�<�cg�(�i0�ĭv!����n�<Y%OU#6}�ȸ���xYP4��B�<`�D7jDlApT�&�iiP�AF�<11/�& ��p��fn�U�t)NX~�S�̇�I�|��}+W�T����aV�F�X��B���`x�#�T���� ��C���Vޢ9�JP��#��E940�	�'�2��	�XQK��67���'j����` ~zL�ذ���z0����'xjr�J3��= �랔#�l���'h��l��n�	���"G ����)�'�?��W�m��X�fJ�N՘d^^�<�S�H)�D�K��Ӯ=<�����X�<�HV	p֐�Wl+J9Θ�r�X�<���z�=x���q���h0BWL�<	��[6k����N�j.|X��S�<���
7/��QpܦPg(=��#Gj�<ԭ��*��g[;C'�ˠ�b�<Aw�B�=R�.�5��4�Ѥ�f�<�A�|
I�$�Ȝ?4���i�<9���&7��є)ڐ�$i�<a��"g���%T�J(�zIc�<��e���r;��k$>�b��g�<��@�� t��E�}�T��Aj�<�R��"0��FL�)2*�xGf
^�'�ў��ʜ�$��-kjƴ�5���$۰م�Y���	�ݫ`戤�'��[l%�ȓ<Q~����[[�p�5K�+@jl��l0tAj��̊_<lت���J�j��ȓfl��@�ɤad��"�Q�{$Na���^0��J�Z f�ȴJ�x�J=��8-Rt�!�q��}���9K$���<����� ���N_� �F��T@ݪ.x�u��"Or��s�Y��]��O�eu�9��"Of���P�1%6$���D�6\��"O��Yr'�3��4�a/�..V9�"O�u��$��8(zMcAo	<+H��ɗ�;4���� 8<T�0\�P:��(�,2D�\ȧ�=�.�0��[�D3�4�uc� %� ����
�z��پk9p�3d� �2�"Op$�jr�j��ba���2�%����"|�'Ô��r��) ��[�&O_�����'K�=;���n^�@�Đ�[����'��`�ى1`�c7�K�K��0��'R���P�X�(Ұ�Y�u4(��s���y��No����v���j���q��ܚ�0<�N>�-O��v!I�o�J�
��yk*�Z�"O4a�5h�	x��Kj@%��z�"O>e�Ӂۏ t�)���ɢ=D8$�"O� � fƠ8�P���կ>C���"O�aw���,�"��J�#7�h�"O:t��H�6MTMЩ��Sx� "O�=�tD��xS��aé�+�kQ�'���:-Ĺ!JL�I@&I`�FB�?�B�ɏK��X�G�O�@���$�P����>Q@/���E�؜'��{q��m�<!�%�z�Hպ�v��Caf�h�<D(R�P-�������6�lT�Uɘ_�<��iN)L��$�C�[?&I��9��W�<A&B���L�i$�ʳ�ȁ��j�<$����HaK��D�� 36��*V�3?Q������ĝ|r�N�3�0�#�9Q���!!���y�̮K��방��5
GK��yr ����1��%hr��'�E��y�`�4j���r�#��x
b��$���y�n�~�Iq��9wJ*�:�䕋�y�v5��)�	�jm�]� � x2��DY�{�(ܓ��!r��q�J�0p�!�AP"ʱ" ��0|Ni�.�9t�!�$�{��	cݠ9�@A�f��)!��.����v�W)=��l��e!���-EMrEj  1$+$�+�Gқl]ax���-�<�RGf
4M�^��B��>�B�ɱi��98��_���x���1!�B��S}�� ��T�]W�ĈE&]$���>)���	b�*x�`L�1�|�3���s�<����MRV��1k�4�A��m�<i���'�8]�0�b|�6dU4G�^C�	1c.<��&�B" XG�c�#<y.O2�} �/��p��� �2�"���q�'u�y���3��Pj����}U2�� F"�y��=�ԁ��R�b�d�G��y�D��N��)�6
{)��\V��T�ȓ �H8xr�Џh� )p�M4n"��ȓ*9�<b��OA6<[C.@,����;m�|#�/V�s2��dJҩE�T1�ȓ* <�`C�Z�@��)�x�i�I>q���	�
$<x5�R�I�fYH��a�S��!�dH�rɦ	��@�%L�t`�ʞL�!�D� {��M�IP���Rs���!��]�M�2Y�CE �UJ�#��2���d���,��TF �7��2AJ�ybg�=�ru
7,�)��!�uk2�x�'�d,���#
Qh���PcA0�X�(���X��I<,*-�F��h��䉳��0�dB�	J! �i��6-��⁅ـ)\fC�)� �������RK=��5Iw"Op
���%s:q���H�a"O�90��Zg�D2sꘈm�
H��"OH���ݨ\C�|+�(Wst�B7"O�hz� �<{��𓰇L
�w"OF��-�+
�@�d�U���۲"O2���	�f�Xm؁7���r�"O��4f�$���0b3���"Of�J�"�?rV�r�ݯ���F"O�@I��{�hS2���Ѐȷ"O�C�n�	7,\�� ��c״X�C"OH��P��w'�
d/	�q΢�"O.���#G0��d���t���@�"Ol�����=�EL�j����������M��pҒh)  ����d-�Q8$-(D�Ha�N�a��ih1�Q
8�A���&D��*"�?~�z%�4�ݴ.�A��8D���eۣ'����L��ȩ��5D��zdJ����� b�Hj��3�O.�M1��#�����0���|���G8b!󲫑�N��8�DJ�sV Fx��'�<̚���2.J�:V$�3�� �'�̽�C�K�g}��E��2��u�
�'�B��E��?Y:�<�T-Z�$�L�

�'�Dy7o-�6��'� �Rx 
�'u��P��������9��P	�'>�ȑÊ�*��}ZF�Q?�8���'����B���8���rBgXm��˞'��}"�'QL$�$�P&�&�H�ҷb�Z�;�'S	�M�8p����N8
G���'#z��#$�7���#�
��9~�!�'Y���.�J �1�4�h2�'��!�bJ&��h�a�УT��U��'�� ���lfNe��̗�w u3�'�|��`^-4'�݋�i8ql�(�O���d�:~�iC�� ��!Z!����)F�'�y��\�GH!��H��z%Y��ׯ%�&q�a�}�!���[[���Z7$���Y��U:m!�D},9J�	��?��+�Fѷo7!�Č�e���f@�5]����Ь�z�a~BY�S��++FQQaPje�@�C�	�s����[(c�I����-��B�I=ҸmG�����r%�TqV�B�		}�4KM̰S8���ǭ?�B�I4:��!�]12���X�HĔ7C�ɄJ���2B�ݬ;��H����B��C�ə_�(0b��/�\P� �i*�B�I�4��	�ul�T���N��]P�B䉶P��CgbIK#4�Ғό��rB䉫TqΌS6��$���%͌s �B�	^��iX�g�b��1���T�HB�	���8X�灄8E�){�-�v��B� ]�P�w�D��<����G�8=R��D����fh�"R(z���K�N�{+?D��A�Ʉ�jzqZ��2hUT�q��!���d��E1��ͅA48"#"��B�ɃloF��@� fC}�S��3ZB�ɖ&�i
��y�LU��AM��C�I�G��P�g߇z� �H� H^B�EdQI�E.=)���`��q�2�	O��HA���;��q@�	�g�8Ջ0c;O�=���,s$Ys �	�%�>I�%��u�<����x:���5�ʪ20�,Z6�m�<� ��7���l=x��o	)}�z��5"O�Xj�yS&] �[B���zW"O �
�H�4j��`�+�s����Q;O���S�Oє��v�`��K6�3W�T�#�'.|M"��D:'����Rc��'�Ry�&�� F��"Q�X� A�
�'�VUBvƘ�N�0�Q�̪d��B
�'����L�N�z�� �/YF�	�'Fʜ@t@$�1�5��*%GD H�'��}��$�9v�ȡl :���O��=E�A�o꼡K�Tu�C�힎�y�M��p�@��C#K�*J�SB�M��y2%'3�Pے��g����
��y��C}k��e��7��d���y�a������&T��ڮ�y�رF`j|��ER1t���
�y�I��pR��܆P�0�RSƍ��yҧ�A�Ḓ�FJ��J)�>�y��/9S���d;8z����H��yRE;c@l����7���hRO��yBe��1غ��d�.O)����y'տ,�h�#(� �>1��$�y��(�N��".��g���r�gX�y�	�T���x�K��`Q� �e�6�yBާ�-x�Q��aʐ��y⯆�<�<�y -ԛF�\�����yr�
	��!PaU�D��!4��,�yĝ�lr�0�J&@��y�N�/�y��'�h�h%	�V ��SM2uʍ��'[T}��ɟI���A狓@#�� �'4�����1�d��'��
�(��'U��C��^L�
D�������'U,͢�MT8l�3$�6�4�"�'�HC���>-l\�i�#u�&���'>����
���M���Kq�vi��O$��D�9		6��dió?A���NЀK�!�dJ��Zx��m5�x@�U6m�!�d����Ć�"�91� $!�I�\�� �5�	6��x1���2�!�$��s'��?�N8B�$9=�!�D��9�X(�	/  ��F�H�!��v?�W�M>`�*U�Q�|�!�D�^����dmF7.�@4@%�t�!�$�}d����SC/����o�?�!�݀r[j���閆dK��pe�%so!�D�N���R�Y]B��۱�Ux�!�D�B���%�e+"M2�&��eܡ��F�E����H�8t���4�y��[���@����������B �y�o o,�y�΂�,�4 �'I��y"E-8%�%+��W�h�`afb�y��Z����IF3��=��h���yrfڦd|1�'G�~�T,�5n��y"��H],�h�"[{<]#��M�y� �
�H�e��`�h�Jh�-�y"���P�b��Z��8{w�Υ�y��'�r4�&`̓7�Bf#�kc�|�
�'�(p
v�E�4��D�C�[��	�'��p�kި5���L�x��|�@�'<�O?牷( `�Ï�?N� 	0`�An�*B�	�X'd�>#y���-@1�B�$� �v���!~����ɘfb�����O@ʓ/qH�#A��ZP��h$`V�KZ��ȓ���I�j�.���2gM�|����S�? $Q���R�0qS!5>��{"O^`��m� B�~�� ��+J���"O��"�ش..졶H�	"<�] �"O$4�Ļ{�6���M�UW:1�"O
�{A?-���C'V��8�O��$[��]ꃪ�J�P�1�i�!�d�
}�y���8�t��F/�T!�d��}^������@����7����!�d��B
$�Y��8{�9�e��Z�!�̵��b+{t���K�!��Tڨ��/E���@�$��=�!�A�6�'0�4���-I\�C�	�_x�*���;౐6%ߌX�XC�I:x(a�W�N�)��1�q��>�,C䉾��(���;L0�]��"�2�C�	�nW�٫!�Ʌ4��%)a�\'Gk(C��
<��S�:[�֘�Dڵl�4C�	^���T��7Q���!���� �C�	�^_:����I���u�DU�<�
C�	+F���ᅭ(�J2�G�G�B�Ie��l(�G��'`^�Yr�T�FC�I%bt	���T�GJEP��EVC�ɣ&l��!��h"daY�희*:�B�	&�TQA�F�8� dC�*یרB�$������N���1$HC�%Z�a�D!
9rD2�*@��7�C�	�ap��9�o[�E9FвaET�/��B�	�N���+ő@�v���%��B䉈o���sR+	1;�~)�"�еu��B䉇?��0
7D��giN5��ASp�\C��-n��0֡�wy.5k"�O$��B�	�&BP@�7DRr�p5Mۓw�B�	7{r\AӯPn��4OŧErdB��'5��Ha�D�v�0D�cNB�	62�De�u���f������՞<�VC�	�-%�i�@lXo�`�h�A�^JC�I%A� ����א(J��%/V<�rB��+~���l 	y��l�EcB�I�04L�d[=H°��$1q�C�	���Y
��QA�PPC#T$B�I1@�aq��ʓQ���T��kf�C䉂7x���@�,d*_0XՖC䉒9� c��J�w,>I�G`H)R�nC�i�#�)�.f�TXp5)ڭ��I�"O���d � e����C�+@��'�vx���ֿ0���	��^�d�ڀ"�'NebE �b�.(����e�'1Z�eш���q%8�T��'Fuh�6W.U��$ү�����'�F����� ���+��W@ȱ�'���H֋�<R��%�2��z3��'Ĳ���H�1J�zAB��	^�-��'	T��{n��@�j_O)
�'�����O�kBμQ�f��PM\�	�'��xk!I��gIhT)�.�)I���(
�'�<�Ul��Fdr"EAh�!
�'f�%�%#K:=@�a�1���	�'����roɇl������G�&����'G� �eē�z䉪� �:K �)�ȓ`�z��g���c+>`��N�3�Rt�ȓ{1B��A "B��,;���ȓ�rx�1&K-8�\	ң�_�Yϊ��!i,	�KC+	ѐq�Q ':��ȓx�D ��O�p��e��H׆A���S�? ���DZ�Y4�9���#]z��"O
���D����2�-O�=��"O�@G�M�7b��zTȁ�A,�q"O0u�����Yk`��p
���"O�	 h�F��q�1�r
�'<�`Z��dSb�Y�b��o���'��@Q�_�`� �B�f�D� �'�Ez���e]P����[�8	��'Vq��&ȊxI�8�ə2g����'�<<��F�~TtP�3d�.cD�'�	���h��Dc�K�1:�	��'�J���,�nL��m�3&/L���'j���E�9��`�MJp����'М�ðjH�2�z`!�$Vq�'�ʴ��LY4)Y m�94����'���!�?@�)���=�*1��'�6}��B���i�wn��Z����'e(��N�S���v�U�Z���b�'h�;�`�|?�C�	N�~I�'b�U:ţӂ?���:҇�3x@q�'���iA�D �F��1��p2,e�'�����@�D�@iq⋉+g٦@��' �DV(��$��0J͹dV��'K�����@���aQZ�$�i	�'HI�p�״Gf�p���Yh��Q�'�r�QI���B|H �$T����'�Dh�Σ~]8l�E�J�F�T���'7�yå�@�q�� $e[(5��+㓯�$�Oh���ܱ\�F|����%)PTY�s"O��m�
�M�w!9+? j�"OpPSbb�=aL�����<k&X��&"O�����N:b����ÏYK�AȀ"O�)Y*X.�,��n�3HI�"O��W(f��@ō+,N�'"OxM�ҥд?�P�3��4r�4�yP�'��	Dy�,�"��	���H���7���y�
Ģ3<�V��=C�64��fM��y �� 0�E�e�,8NAQ(�(�y��R�|��j�:����D��yB��'}����
Ƿ3���UY��y��
�L�P��g��Aȶ0� �!�y�J�f������ ;gnZ�o��0>a���?��f,p�q�I߰{���c�c��x���(iA�.}T�����0&�]�ȓ./Ȩ���"R��ܪ5J��]��y�ȓm�р�	�C���"s'W>�r��ʓF��=��˹<<i��e��B�ɥk��a� T	|�j���ą�uB�I1uGP㦢�'rjd�B�kV+�C������'H/cqN� D�\i���/OD�=@�=GN8T�e���yq���$(�_�<9@D̈58"9x2�ִzMKq"�a�<IT��6
���qF��1�,{
�E�<��4-=ެ��ғ^���u�"�y")Rc� =R�,�Ce�	x ���y҃�0dO�j|��q/��|������?Yg�Ju�����&�`�{O_~��)�'N. <���H#q*�٣��/ެ�ȓ{��Ű&�B�2�*
�
ݴY\�!��8N�B��3sn�9rGa[2Y��)�ȓ|�b$)�f��y�oS,
���PL|���!���G&I���K�<�R��q��"��\��Nt���}�<a5g
�aP)[wj�2�|œEx�<� �A�[�.�H�h2� Y�.���"O�i��i�?�ҵ��&�#'�Bx��"O\i׏U.p!Q�ۨ��Z"O�qQ'b�4�p���>��!��"O�X��L�E2l2�#�R&"O��	"+��>f�`�M��}v��˃O��$ӹwT0�Xv"׶�����B�7n!�`ަ���ɶ0M��S"�!��:�`)`�@�n9��nW$�!�E�I��Q�n5��MR�^�!�׎i*�u2�e	�]-�;�7$�!�� N��1�^� �Q-��	=�1��'� PZq��Z}f��`m��H�J�'B�q���$ra�P:�Cv[�BO`U�$�߉tfA@���`��9��"O��h��,[�~ �U�%�\a�"O�JW"�jy�͉�υ)�p!�"O����C�lɸ$�����m�2"O衋Do�)��q������"O\@(t�� g��<@`Աz|&��v"OX� �
T�N���a�b��8�:O���$�??�8Ƈ	 T	���&��:�!��V�4	Դp�Jҏ{����RD�
�!�dC\�~��5�ǻk���p6�݋`�!���M9��:vNI*�9��<t�!���$Z.h(֦�Q���#��!���5�sƆY�]M
�X�Z�Q!�dʏB|;���mb@�&�ǆ?%!�č�W0�s��	�HwfE�Ʉ7u!�D�(@[դ��@��!�&S!�!�$]�5[���5!���B�%��iM!�ĕZ2� ��2��a��-
6!�$62~:D*El�'y{Ҝ5l9'!�ĀR��\S���c�����8 !�DU�QS�5�Gd��%��Ƞ5�18!�ė�v��p٧�R��,�xw�T�~6!�18�J)Aw#�f�rQZ�� r�!��L�aк!jRl��Z����!v�!��V�|�ZG������C%�!��
�ؙ1��P���*@�%X�!��E�G���j`�#q��q�*{�!�䔚��˗[�Xk ᫴K�!
�!�$K�~oĐ���ѺWm:����Y�-�!�F'Z�r�@�~6���K�!�$­'w&�� ���<E��@t�ۈY�!�Ā�k������	=vP��l(]E!��щj��C��|����+��YH!�$��'^�ˠ���~������%"8!����j�
�#'�1��*�](!�LK4d��	��	tDyq4�X"4!�D��\6 p�PJX�4�si\�n!��b|D��L"1c> ��"�K�!�D�#�zY����Ne� �a�!��ȴ@���� �#\��0	��ɋrp!��28v�2熀�c������2x�!��]>-]���2�P�=~��Z�N�)�!�D]�z<Zp���Ǫ'T �j'��.t�!���1!ZD,�FN�l�ʔA�!�{�p�$F�R���H�[�!�X�{WԠ���b���QGÒ!���{�(y��V����Յ�|�!���
9RU:@�A�0�d����لȓ
��d�N4�i͓�؄�pY�Y!�-�j��錧jD�ń�S�? ��3��4^R¸zG���d�"OH|is#�=S @��ۭ (�ܲ "O�"�e��i��順@ץp���"O |A&"�+ �_8�I�#֭�y�77�01�١U"\�g��yR��O�p�v��H��E!Ў� �yR�ϻ(��=��a�S5<�قj
�yrD�~^��$�Kd�2�d4�y�R�:B*e!e�E3L�&�c�=�yB�ٳy���{���,D$Z�a���y2B�cl��w��,ݔ,��JQ	�yB��':��aT7+Jk�Ŏ�yB���|k�� G��Ra��#�MH��yң�"uD�zbϨL��IS�g�/�y��:٤���阿GJԜ!W@���y��!Z����c��,>�Z�Yqg��y�*S+sPᘷ�U!9&���h0�yr�
�P�*��%��,�B�%lN��yR� ��")�881�����y.�c�r�����N>�T`�E�y���E�R̩d
��M���Sc�y�ƞ�9�<XS$��
8�>�+� \3�yc��-M,)�Ōy\>5" �R<�y	�`���e� 9j}����U*�y��)k��C�̂"Nɜ�h�K��yb�ҕe6UH�̓p9��Zd)١�y���Q�Vp����8_.<`�3i���yO�tCN�����*��D�y+ŵ���"�,�xU�ʬ�yҊ�$$��`&T? �,��3����y����Ҽ8Q���s��;���y�@ !p��� �mr�ظ��;�y�F��wzx�S`JLc�J@2oP �yb��o�1���B<[�ۡ�C�y� ����x� ��P�d ���,�y��]>r�V%���C
��σ��ybI�!-���9�H�:����-�;�y�D&�@5Q�C�?8�p:���+�y�M�Z@��W��-�QN�4�yrjQSp�iE�ҏ+��\�k^	�y�G0x�r�@�i�5(^����DP��y��W�@=�s�X�&��T�1����y"��{�l���������y�̀ ~*l`!H��T9Cgԭ�y��(p喔 ��"�T��R�yb�E�yp���H���e%���y뙂1�Ƞ*�ȟ�A�$��%�6�y���X5^�����3f�萣�%]��y��+���;ŋ�XB�2�fԬ�yR�� B8 �i\�I��d v�[>�yJ@]����I��>@i��Ǘ��yB��\�*L��O�:*`(b�U��yr�%E���^���0OFw,��ȓ
t�U��"�ȹzW�S�<�����E�L���DD��r'��\q�'���z��K�dېɛd���v �(�'�� ��7x�x@t��4J�L"�'�PX1�+^�6�Dy@���'?��C	�'�|BǡW�#X�)c�۳.��͊�'{���A����
�M�o���q�'�x̢Uz�� rG\���'c6�A��D�>P��b�(�)�!j�'� �q+޹wi�,#�W�x��l��'B���0� ��ZE�
q�֨��� �T¢˂�!��	पG�K¾m��"O��#,�=�"msIO�Rr��"ONȪ��"�p=��bA�IΡS�"O�(�E��*��,��#�?[b��"O��'�-���"�.f��0�"Oh�!������!џUnj1�1"O���5f��_Y�HC�֛Y̸(� "OttqU"�y�T�pcֈ���S"Ov��v�E>��� VC:t!��"O �A�/�\<,���`��=*�)+�"O�Ͳ��B�/�(��H�8S:�C�"O619s�!�(`h��EGl�"O�|��c�Z�Kd� -2�#"O �J���$|:�u*ਝ�)0�%�t"O �AO��Dd�!	E3,���"O�p�k��|�P��t�L��R�"OR��W>�V$9G��!c��I	�"O4ݪP���i�b8qWB]��*-c�"Ovr���&���p�͸A�*Z�"O�!�ê�%�{w7+ؕ �"Ol��b�/y���"�քlv�r�"O|�O��?eXQY�.7QQG"O��ZR�]�S��Cj�G�MZs"O�,qV�6<�.��U	�;��8%"O�m�0��rce`ҧ��`iL���"O��4CэVL< ��P�eU���"O H�цo*���冺;8�tb�"O2(�"�7u�l)kF�_6y��Xp�"OЈ�3�$@Q��iw�45-�Q�"O�|�E���|���]�F�8�!Q"O"�VgO!����R�w���"OD�T�������'Š#�|�P�"O��q����t4��\0hp$pj�"ON��G�^�j�f� fG�*��Ղ�"OD�W [�]eJ	"�n=\�J]hf"OXX��R݊��bM�	y�4t9�"O,p�7�'3�V����]0��1��"Oi�rJ� G�E�0��ŃWnS��ybn4Ö�$ł�	��:�%���y���P�!``˲ٔ�;pD��y�.\;]r!R���X"��.�y�e'h��Ѧ?���p����y�ߜ9����b��6j�h�A��y�f߫'5�yMG�3�p��wȌ�y/�5�:�f�ư%=������yfȴ"c���"����b�'�y�.^�ΒA�,��D��8�����yBNjKDZyW�B�dT���2���yb���-Wl�:&��*�̓�Jˣ�y��ğ"��s&�-7� !�����yr�I�3����t�Ӏ��k�J��y��f?JIU`�;����ybb�/q~��ɋ?xT%�P�7�y��+t��T�����m`,)5(R�y򍇌վ݂��\��-˄��y�&S����,�S���%��yB�6��  	,@���z��ܑ�yR:��m{b�O
a���)�oB�y���2_�0Ъ��C;�=�r�5�y�Ä5�"�g�2h�x<ysN��y�h�!Us�8:f'�[�.0�#���y�	.X� �:�
U�2�ӱ��yG�;������7Y�hJ�	�y�lYK�Xw͝�#��L�4l�6�y
� �liT��*jƼz��K�8���a�"OL�k��Ԃ��}���Oyb��'"OX�"+]�)N �T��K�L�+"Ov`�@m^�JMb� �ێO��LP6"O���0��0'h�!��1;�m1�"O�p*aǎĺ��3g(Z)F"O e���� %��La#�b����"O��#�u�����%�EyU"O�ҥ 	  � �pjÍSݸ��C"O�`����3P��Q�ĘMz�1"O�B�l7_瞽Beg�%m`8-�`"Oj���ř+�$���@�E�"���"O�Y �
�<�H4B��E��Q"OʹUE�u�2@�QoO,c0p�u"O�R��N�s傥�TΒ�����T"O��2`���/�@@�7Ύ�{���r"O*%��Y�J��{��ò�Fɰ�"OV@B�LF9\8�qGnM�" ��"O�ؐ��r\�8�bl����jq"O��AB�%�����ܰ(��g"O�z�`�25��x�᫓j��tir"O�����[�rQ�'�*i��cq"O:m�G,W7:��C��?,��s�"OBu��E'\�T-�R�L�>0�	��"O�)�BS ^	4�5v�:�"O\$��&���6��끿|�ꭂ�"O�q����]E^4��i�3e���1"O�	s'[�6|�D
4'ɓʒubP"O�آ�eR�?:�y��V�Z�T)�F"O��a�Z�_�|(�L��b����"Oʡ[�*����E�]0R"ON�8�!U(Eޮ�j��7I����"O�s��ޖ-�<	��`�$F��#E"O���d��
{��P�-5�nQ��"O���SN:D�*)�O��DiH�e"O��"D�<1q�P/��nzJ004"O>��ʞ��.,;�M��)v��0�"O�� ��2T^�	�f��as���%"O�A�uc�4���OD�2m����"Ot�P�F�z.�(R��>KJI��"O���舋ø��mY�fE桋�"Ov��D��a�E��LQ�b(��"�"O����΀1&P��Ƅٷq�=ɶ"O�Գ&���V䤕���*�cs"OR)�$㋈X����ь�v\l�"O||!NDA����(�.$��2"ODy�dȐ_^�z�N����"O�آ��� ��Q�\,h�-ka"O�����M�>��І��ڰ�"O\a��
���KR%��
]��"O����j��'Ŗ+:�Y�1"OH�S$M�t��8�b�^=�l4
�"O�Mr%�>Y�$H�EA���$Y��"O���d����<8v��[�A�"O�eK5�C4D��P��k�������"O�]S��4%|l16���
��"O��c��0��CW�Y�c� ��"O�A�ԈW� v���5(VհqbA"OV}K'�2!l��3�D4�@��"O�	�v�	@:
U)G�òF ���U"O6u�aK@<$[��#�FF+��A��"O����k�Kdp=����u���i"O�(� A�T���A`��[�4�S%"O1�ဤ3�L�/A�6�4L�6"O� ��iG�Nx�3�[�\��C"O��ct�L�����M��1"O�-q��H�,���2�D�ލД"O~I�"	ޔ�R�Y$��$���bC"O��Jׯ�k��������"OFձQmۤi�AT��5�"O
PC�H�/
��2FD+I�89��"OH����QװA�`ǈ��X��1D�ɕ�͹#�<z�/�^�HQ�K3D�|B��3�e�rm��>�bD�6D���F� 1g;J��*ܾ=b�X��6D�"ҋ��CD�dy��\�  C4D�H@�-�6;�jlo�� ��a��
�c�<Q`D� ����%���	�g�<qmQ8mTr��P�%&,-p�*II�<�E���0�慸����#�CG�<!3��P+v��Ï��������@�<�#��>ZiPC�o��D@��/q�<��O۾lq��VNӝ9�p�iP�Ep�<�1��N����C� *�Y���u�<�A���c�v�ҳ�Ǻ=>�9��]�<��L	8F2p%����a�1Sm�<�䋊#Tn-�p�4{E� �Β_쓭p=9%-�|� =�B�̼R��\�W"Hf�<�	_��U !	ߴx����e^c�<��L�4�h�
g⚱VXY�BF����>�,V/��"FI
�g"ص2CNU�<!��T (ӄ�0o[[�LɃ'�~�Rё�����!H��'~����#�,+���@4"O\I��߆.��a��6n�&Š�"O`��V5 ����G�D�t(w"O�4��D���(�2�ǝ-�i��O����� �0�q#S�G:�����
�!��$�^1x��ʛW7���h!�D�SA{'>ej��R*S�!��&^0�@�m�0Ơɡ�5�!���L�訪���7��[a���!�� �.8�!o��B%�6k�>u�!�Q�s"x� �`� ]���A韻<�!�Ę �\����>T���s�ɰ>?a~�V��+u��|ϴ�ї%!$���:�";D� �`
^��acD��Xd��{c�:ғ
6a�DE�~j ��e�t1�FѦ�y�E� "E�tsr�ΜV"�۲AC��M+�'M�O?7Mѵl��s�#L�z���j�%��b!�_?w�ݻpk�l�!�O
�';����ɾa?|��$�+O�\t�F�ޮS����D����4g���˴lڰS�ѫ��_;,����ȓa>����@ьBdy���Y��mG{��O� ��BAZ��(Rf4R��!�'�ʜ�aΓ�c̭y"��& 6-AM<y���	_%cR�8�4*@d&Z|!$���!�$Ϫb�:��d�K�a��z�d	�p�qO��p	�"gH�)G��'y.@ٓs��@����ȓt�<iBlCl0j���E� E���ȓ<&$�v,�����MV�>���ȓ2���c��:t�E3�.'~D��9ϐ�ga��<c�K@�E�n��ȓ*ʘt(P-H��l�c4�K3x��ȓL�d)��đ	A�|�4��;t�G{R�'�N��.W$a�Rݠ���-(��C�'��PgZ�!�����4�,�J��M[	�O��!
�?Qv�(�aj²%� q�ȓ4�$|w& !��PY���)�p��S�? ����n�L��RU�`;��;�"OH�(���H��� ���hKe"O`�(�Bȯ <��BTO�r`�%�Q"O�F� `<�k���jk�Y�"O��EF�7K#F)X mԿGW�-�#"O��r�\��;lͅaE<�!�"O��;�HD:�B�"���"O��(�KRFi�dJ^e�#"O��c#ÃD%�Y�##�%8"O�l
���a�8���@>}H�@F"O�1)�.ζn>� Ќ�2bH�x"O$����&6�
�K�
S���t"O��Z0I)��K��2�VD`�"O�9$�L�u���
��	,�4D�"O�4�� �~�ur�(S�j���u"O��M֭	�� �ȍ&B]H�g"OxEW�P�t,���Hv,��"O~�����+&��,
#Ҭ23`x��"O��KB�木k���l�h�"O��`��L)�X�U��z��!��"O�1"Ri�.��� ��?��B"Oƌ�D��Bf�{�셂$Z
��4"O�壤�¯.�����H DFy�7"O,ܛ����
=����:2���"O��;�H$�N�� .ek~� "O�����ζQ$�P%iW���)y"O����gB9<�Q�7'M��D�i�"O���g��Ƶ��y�x �"O�1:�,	!M�C��� ���D"Ov�����j}�U��5m�����"O��� o�g�t7���e6��"O.���G�QC����	c�9�"Op13���v�X�����MT���A"O6���+;�@�S�Ŵj�t���"O��ч���X���ǖ>vf.�3t"OBMH�)6FW5�"������yB�ɏ*�PУ��)h}K7$B��y� ��j��Ĺ$$�	T�4���D��y��)d����m����C��yrmh+u���	9�y����yRL�;D��pu��4&|���8�y�k�#\���df�7#�FC�
]��y� 5uX� #jK &j���!IǦ�y�X/��
v���#N�� ��y��0e�L���cH>-3d��,K�y���T`b��D�.).ތӲk�9�y����pƴͲ�) �&�Ȃ�P$�y فRw��D���(>��S"���y�mJ8�I��A�o��d�1�y�ׇT����_d��cF��y�e�!�P�:�cp8�3N��y"ŗ����:�f�\�3��y2��:�2�Jc�X�+������S��yR��kCf]jt�Z�<,� r,���yB�7�`��pi���m�b:�y�#�8��B��?r�����y�K�#��x��E� ̆�y.ɦ]b��n+옣�㉤�yrc�(qO*�A��d�x�Y�Y�y2�Y����8`�[M!Toӿ�y���s��d�E�T���X�/Ȓ�y2�>��;VFRX�+�区�y���%k��D�Sl�/h�ͣ$S?�y2��6��i�Ā��®)��lX��y
� I
��O!=���p��	�B�f"O��K5ҙi���� D��i�6"Od4	�Ђ|<n����ٌ(1��S�"O���A+Tv�D���H�$���D"O���D�x�2�����:8�.]�3"O�L�Fi��)%�X��H��Zp����"O��gG�cB����2�6���"OnP3��Kj���$���� R"O�
pΑ�W ���?�
��1"O|ȹ��T�&�<�&�G�j�(�"O�*T�O�
@Z�s���C�BR"O>u�`�
LD���NY�G�l��"O�86,��"Q���I*��u��"O�z6�A����+l�X�"O,a��5Y�zE�eNW�N��!�1"O|%�����Y�R8ᣭS����R"OV�0���lzr��%� W�DQ@"OX��2K�&1�bV�`�E;"O��� �[�q�V�B���� "Oejt��D���b!A�t�h� "O��Q��2sd�L����(V�|�"O>xB��Mr�͉m�+�"Oz�D�
�2"���&�K
j0�@`"OIÃ�֩'sB!d��A�(�1"O�$� �]��n԰D�d�"On�۔H_5	~���[a�^���"O�	 ���<d�؍�� �<!tЌ؁"O-aөM7�8���.E 7f�l�@"ONM��l��|�tu(�΍�}��l��"O��&�2��� ����
bIk�"OB��f��]V��b�u����"O�<�
J!�U�FK��4�"O<�EE�;� �s�ڹD�X�;!"O��h�P�\�1*�,�d���"OQ^(��Ucݯs�z�x`�ֶE���r���Qo�=mH���o�6�=D��؆�5F���%�"I6��bӮ<D�Hr E�c��z3!q�Tp�y��'V�	>9�F��[2|�0���E�*�9�6D��Hb�_)e�숻�A�?3x��M0?i�O�����Ɯ�F�+8܀��Bğ'ua~]����+�QG��rJZ;����D.?��gTb��lI�`�u�X&����vy�L\��ڢ��.3JJ�K����O*"�#E�e�4t�qg�0`ȥ)�#l?A���~�N�t��Y#�M����Z��jeH7D�S�h��h?&�[sΏ39�:��5D�|)����
�a�·L��+����If}b��#J �s�ך*V$�B�gG��p>O<90#3=��χ�:�������m�'�?��Qk�!(���K�(�s�4D��
�m�h-��K&BD�)����S&7D��au��5T��(�%PK=$��(�O|C�I�J5�{G	tP��/�#s�����#�I+km��a�
G�hھ�+g�;'�C�	�B�LՒe��2/��(��|t���<�M�d��b׬���7q��!%D��k��фO�"ESį�,h���m-�d2�S�'a�4lKRF$f�="�n�?A�,9�ē۔�R��.0b��H�P�f8��"O��C��S�,bXa���S��cv�>Y����O�O�5̒'^<��{R#ȤY�TT�"O���	2mVx�rC��>�Y��i�ў��.�Y*du��[G93���*HtD��S�? \�*�Vq��p��֞0,T�r&�'K:���	48�T�*i�7Hp�nݷ<eੂ���'xy�R �.RC<��*	4�@@�'�:d���S��h����ׂz�'�
9��_�
$:A
��	����'a��y��F0ղ՛A�S�L��5q�'uJ�i���c��5���Q�Dz���'h蚱�>V���+c�� '��Dj&
.��ȟt Z�,����u�����'��� S�*Fi�^%�u`���T��.D��Ҁ��6H�B��W�F�p��`bF.D����Y�AK\�pː�Gז�rPB,D�����U�>�%Y��>}�4:eO/D�LK�A�9Y<�yPC��{Ԩ��w�,D�t�0�	Q�40GFM+\,z(�D D���Rh�Qg�th� ��b\�,צ0�O$"��w����Ń�,����Ð�g�0����<)�U�,�T��f�a�clS# T�G~��ӻ*n���lD+7�\��q���xC�I8\k�`�R)U!'�x ��. ���I+�qO��&���U���(բ#��X�l
P�<Q��N�K̉�j�.�[�L�<��O$��L<��M'?�a�dФl�"I�qj݃{N�3�h$LO�7q���Ol����i'��1�n��0c&k��4�S��yr��F:�/�i����B)ү��O��x�O�$��j[�=;����C� -r*yß'��BgM�D[$�u[��ā-���yr�'M�O?����No�(�JV�T�Ф��@<D��e���q�d��0��eC\Z��;�$"�S�'A��9j�$[0a@
�`G��M��(�tx�B5d>���0�߷�,��?Y�P0hl��a��
S�KA��:����ȓ$	ԝpG�T���ʄ!	�o60���vC�M1���Q��x�����������/6��S�OJ�����|�F�`&�&U&F<0
�'!*-`e�L����!;�('���'8h��#.(8`��؊@���A���:O�ab�O���� �r��H�*�veK�"OD�R��� �,�ɇ�i�Ni�"O�I��ƗrȖ�kF疎6P��2�"O�(��H��6B�� ��UB:T��i��IO���OU�p�Τ:�3d�ȯ�r�)�'� �
��B �H�#i֥��{2�'ߖT���0s�,��a�J��}b�)�	��p�J�y�'��I��`rT�Ԩ*!�dE�P��d)�iy>��ȑE�t!�d�;+��P�K�9	:f�+�oL�|!���x�fL	'׺P�py���P!�$�p��!M�#t�Q�/õ*M!���"c�X�AK�j��3U�@��!��L<i�=P��h�2���!��_8�i!����%�L�i���H�!�dT O��Q�/Q_[<�H�e]2j!���q�j� ր��5l�Ӈ�eU!�$�.q��P�$H�1ub�� �!��"A����b �\0�)J�!�G1Z}HDBg�1(��e�#]�!��86ġ��$"3��x�ޑ}�!�$l�uiJ?N���ӈƮq�!�D�dyt���AWEŸ�2GD6	��y���<m᪔  	�v�b�#͞H��C�I����I��9;��0BJ�+��C䉤W��8���J%~�p"�;n��C�	1~۔`Q�땾@�����X�i�6�	æUFx��)� ��� ��M���X������$�"O�ґdE�RHRs&�}k4�┟���ɰ)B8,CD��-<���q�i�@�fB��! ��y"kB��M�Ǝ<�dB��~�!b�ش�ȍR��>h&B�I�M�+F��Rڐ!�.��9�����'�f��SeJ�����=3B���,�O<����$2��sqGĄ&㺨	�e��D{azgHT��'M������O%�:�p�#v!�D�P\xy���M�=��9	��_�TXqO ��V�I���Ɇ�tQ�8�6%�T��K��M�L:��duG"�ᵫI +8<�s��̓X�"=a�X��${$*G�Kv���`َ�x�ȓ?BTK,R�U"�5�cjZa����ȓ{����� D��@.�|<`������Վ�/G��2Q�D?b�܄�L�I���U��Ƞ
Ĩ��]ɸ\���]�O�������=\�Iꠊ7�깅ȓ�,y�ύ�/O\!z�ŻYZ\Q�yb�l���Q�6L�p�]�:�`M�1h
6W�.P��A�B��\i�%��4.��1�T��\Fx��U8�x)4e[
���7�	���E{��1D�ؓ!a�M�*��4��z��2�"D��9�٫^���I��$�s�N!Ov�=iu.�V���[�h��Y�p�Q��G�<Q��П*v�*#���)�D-���l~��)§��Q$O�3z@�@���W20�ȓ,��ٱ��ՀQK2���CUT��M�ȓl�i���v��
ە*,�ȓt���#��pp^H��Bԝ�P�ȓ}J���C�e�ʹ�@���fl�ȓe�:�8�E� =>� g	
 �J��ȓQ��X6gB,,�<<Hw@�8!M8���|�1뇖+���+��÷c�l�ȓd�"�9�	l�`��L��JI��p���t
)�<3"45�����r�2�1���j�(��J��t�5��x�<`h282�A%�o�x�G�o�<i��EI�h��/W�`��R�@�<���_a���x�뇸x�����H�<A�'�i��t��3-�X�M�I�<�w*�:$��-��@��&�~� �Z�<i�Kx˺�[7L�*+�0 ��|�<A����<�ӵJ�$��sEGz�<�%�?a��@�u�=������s�<!4BQ0+�Lc�J�C�vX�p��p�<)S�	&��d�f@8ahȓB�0T�� �A��_��A8��D�1��Y�&�6D����N�N�ܐ򢂿b)ly��/D�\keI�l|Ҷ/�#>)\ ֊*D�xF䔌MX��(6�/	���ZG(D��"�A:�}E���J�nY9��$D��a���4��m��FZ4&�=xP� D�,h$���6Ԃ�a��\�)�����!D�����aKXq0�'ڂ,�ո�B4D��Ʌ+1{L�r��ʤKs���UI0D�@��ǉ�);~Q�#�[� ;���F 0D��cP9�1��Lڣ k��h%�.D�@���FT����-�\v����D*D��b��={��ԡ#j��-�d8��n)ʓ~ሰ�)�|����ӊJ3*�z�'<��R��}�X[r%C��5��'���i�OY#����d�9A^i�'�8�A��)\��-R!@���T��'ؾ�Dư9X��Á�ׁ}��S��� hS6&ɂ���[C��2���"Oq7�J5 ~�@'e��fˢ1�"Oa���Q$�Z	�"&Bm�Vei%"O��s����dL����ZXz@P"O�,��!q��5G��	6���U"OTIcB��
'f�t�)Ԗzj�	�q"OzLz� ��:he��Y�pX"у�"O�x�!�A9gh]#��� YP��"Ov`C��G dy�r��3MOL���"O$eC��I%HTV�TNˁ_+�d�4"O���t��3Aî���^ϼ���"OLp'�@D��,�`��W� ��"O\���x>�ۂ��:m�vmQ�"O�Q�F��*q�� `^�S�ڀؒ"O�1��ЧUc��1� ΃k˨���"OBpp腓$���K��(x�@5�"O�1�U˖�a�tŁ��S2Ef��T"O��5�K�ECC���`2���"O�}���%k�6��rL��B*6(�"O����ӊFg�ap���#��"!"O�uӃK]��.��&j)+���)0"O\��F���{FDM@b��!"O��B�@->�НD��Qj& :1"Oz)s�4�4@4�(�(��"Or峑m�]by2�	�#H�Z�� "Oz5��E�D"Z���.~�,���&v��I�o0]>X�I�O]��ȓ!d�P��Lm�)�6��"pVr�ȓkG�Ȉ���R ���B� �مȓ�*������z��;�'ۜI�Ȕ��D��	7�O�q�@hC�f�	�α��1��8Z� �:
\Ru�f�ŕ
ӈ��ȓ`�>�B$�S�/��	�$��.@y�PFy�狥a�:�F�� �LG(b�l�6l�R(��%�:�y�Gq�dmK��H�^�:yP���V~ 8��ַu�ɧ���D�[��#%��d���ؿ�!�$ʚM���KP����,\6"5�-Sgv́T�
K؞D:�b��V��E:c̉o�R� �$#|OȶjeF>T*۴\s��*'�'�B�JV�V5��� 5�EO�-p�{�[�^�f$�?��k\�br�AU�>�'Q�d�!#B,g��1ip�K^���ȓ<�@��^�:i@��׋f��d���s̨�}��h����!P�N�&H�tf��v�;l�!���*_(qx�Mv�V`*�@L�'��'҆�l�0�˅f؞����� �lZ���B��is� /|O�$�_51 ���4*&�X�'��S����3�W�#�P�ȓ`(I뷂O�%_��8eF��: ��?�'��=	�x��/%ҧ1�N\ڇ�
�ޑV�#ej���j�R��Wd�� v�| Q�	1Ĝ��*9yO�P+B�>)���O��@b b�p!�"�bX�Q�q"O��ڇ�
�=�^ s��%
�Ա���'٬���3DkD\��I�R����� �.��b$�]rw���Đ#kꈄ�s�O��a��
U��Ӱ� &/��	t"O ��4��(ff��\�Pupv�	fe (��u��HS�.�d�v �G�� -�B�I�r�Y�̀34,��[V{bB�=h���qOI-k�0���✈^lB�Ily��i�+H��@�lΡQ#`B�I�k�Ĉ��\�Y���$�I-�TB�	�GȰd�c/Õ&���h��#�j�Lf�ɹ~!�#|�'h8��$��rC�f*���'ۆ8@��]��}#��L�;A�1�&"���t%�+�wX�����
�I�~�#���9ZuP��#,Ox�Pw�̨\|�ƫ�Đ�ۇ�b�!��^�ݒ%-D�� ⠀G#U�r��F>���C!�x���$v��'B��Q?�Y�
A6@ R�� bX d�H�q+'D��2tc_�/�F��e�w7*�	�.�+E;��[�Ԁf�����_���ƱyX��/?��bO�����
�)�������R���Fb��������:Yz��$W>?~�Ƨ" u0c҆��!�ay2,�.A�< �� 1A��ײO�Br��!Vk�	+%��j�!�P�s0�X�/�::���� ��<ˉ'v��a�A�2r����=Bm:!���&Ju�I�O7��C�ɦ�I�����jS�����J1(�nq��a�5j���+*��`���L<!�&�/U:��B������lBh<��ဓY�����̎-��tΖ*
(�u��Z>��s�PY�0`)�g���B����k'��N�����	
sN��g}�K�.��@�cN�OѴ4yg�r9��J�)N	8a~�K�R�q_��9EK]���P�	˓:�h4�j;h��J,� ��ѥ3�R�2vH?	1���3�~���gK%s^�B�L�'x �&����F&J�P E�ӥ *�����̺C�&�+E�U.G�B�u'�ś@��x�����R�e%�'�]�U.����n��I�,E�%�J����DÕV�H���w �Y1ȝ<��y��ޏr*�Ia(}}�p�U�8��ig-�M=v(�e�Z\��\�vܜ���	P[dg�V��b���Zp*�%�0��̇*��@:���(c�섩�jP�X�d�2a[>�yA�M�m>���>a.f�,D���ӊ�xK��;a� �N�#ό�9����K�t�Q/�9"����}�7��}l��=��U@7��;voTq��j��hV���
A���1(B���т�C7r��V���6x����.��!$��h��%��퉠U��<+�͗�J�| !���,-�p����	l��}B���}�hui�p��T�bT�����c+G3w�`�=/Lah�M=�OZmH�K0���@"Q�f݄�b���$#w ��K��9K����e͓rL,�Ĝ~2��/�!�R�� _��%aAG�<Aqc	s'Ѕ��A�6��U2RŌ?�� '���^�*Z�"Y�4$?=pӊ$ ]�0�,���)��O�o�	[DGN�<E��ɔ-��ܩt�<&�"Ȓ��%'� i���Ji�;b
��:�V@j,�d*>e��>�hO0�q���zkb1�(�!L�4�A��;m��c��ؕA  m��A6�a�bR&G�xa��b�;+<��q �Y5*E"���:+R��dțo��ZvE��Icb��i��@,��2*UZ��וNg�)2��L6=@b%��ѧ7�zm��V>�:4�E((&�2�K)E<i�FE#D���� �,��E@c��Z��d���j�T��)^�5U���Unηtޱ���|a+�i	�ϻ7�@����5���$OX�ttĆ�ɘ7��4?O�Z#�
s����D9d�n�pLU�R�$����P��V!	�P��ɓ"v������ɽ��%ZBb�`���F1�'���V��c	!�2FL�u�T��j���h���z<Y� G8wg���!���Mj��� �	x �3&�mx�`P��\ ~�rA����3 骅ʕ���7�.J�����A&X�H�� �ѸB��Ɋ
a\�%�U꼻�"Ȯ?�%yVHÜ&䨱q���h(<QQ�/e��@�D
'��Ku�5x7�|�R摍�@�`⨀=TD�d��#*o�� �d�="@�U�<�����'٬\����qsු|a�dv8�49�C9h脓��'ڴI�r関.w*m��A�Y�X� O|d���ShJD���̦�٣�,ATQ�����@�P� [��A�'}d��%�MK�^ϟ��� iD@K�"-������t�lJ�`�(!
e
U�(($���"O���dI ����T�Y�i�)(��H���Ja�u��[�'��Ti<�b��7)B�]8�̈��D��5dn�8BS	�(B�T`ZP�MǃCT�)�ꂓ{����� Ći�l( DE�O,0�珝<k��6	YY����L��s�#�#45�9`&-���p<qVnIO���PǠ����c�)J�ұb�V�
�`�kJ7&p�b���*(��c��'�vu�F�
�.���M4 }�lzL<i�GۑjE�T��Ob��"O� ӄ��������	�+">��s�X a�L�*O"���]���8��G�\@�٥2���\C�����K�"��ğ�Aky�LZ��4��K�=1�!��$E���#F*�+z�И2D�4i!�$ȇZI>��TB	4���`��̶9m!��D�b�y3���ˆoN�@�!��a�\����D(ӂMb@�v�!�_x-�P�O.\�rJ�Ō ^5!�]�6(�����,��PvD�I!�� T���"֎s����
�*#�>9��"O�*�!��)�}�tK�/e��@�C"O�Uh�JO�G��j�+s��ӄ"O�D�L7�@`J�:j�x�>O�a�aЉ�p>yuk�,[��p*�&o��uB&�w��h�k�f�|�o���SnKm����F,2����<@8�r'���E�I�
�!�c��R(�	vM��@��8<p��AMJ��Jࡵ��"
i����"j��ɖq�����<I l�g�c�puY+Y;J+���O6�F��O�qcw��,v�~8��/4r�p4Y4�I"S�������p!�����H�4T;���f��6�DP5�$se)F����jO]H�q�
� _�ypf|�D�9è�����U���@,F��?!�eh�6���ڳ6Ф �wB�<�"FI.>8�<�d��v!�Ņq}�A�'`:�!��)+��IAӄ�ߟ�j"�úA�~�ɹ1���87K*i*Ɇ�I�W�|�������P)���T� I�R�� 00�I�b�ܦedi�!�b	D�4k`�Ē4G����ę<%aC�?�#�lU�UO:ڧT?t�H��!-��g,̝?x0p��W�,� �b�-~����c�º۵�!�L�$x����bT,� D�j����	�I/�(�?�O(P(�ڨb�A�l��0�cE݈gX ��7�^ԡ��19P܅��I�:�c�nV�	pl���P�J��"<�qi��� ��-O��Bt�����ƞI�T�h��T�D���"g!��1����#�0@�uS$GG�>`�'�(��f���zʨF����{��Ѣ��Y�����y�I=kCƬI��I	����KօH�@̛�>9g������'#0d�CC�Ũ���������{�'NA���T�<j6�#%�D6��g`��]�^݈���zx�0��D�}h2�C'A�c$�%�'j),O�l0g�u�BxC*O:Xɀ�D�y|��v�W�Pa�(�"O��)�n��V1��SY��ؚ3偹�䓁Ek�+ȁ��ө&ߒ��0�	 a�u-e�Լ�"O�Mr�L/.�H��WN�5U�@<,X�Ez�{�A����)�f����N�
���)5%\�C��S���(�I�#6�����I��C�ɧ=iN@S�+�I���Q���C�ɇp�2��f	ɶ=�֜���[�f��C�3��Hѫ�%=��hgeZ#g��C�ɴe����ϝh�%�3�ڼ)�pB�I8S�����J��io���1�Z���C䉍+�툱*�*/�����g�%8dC�ɝ{ۼ�E�W�[ލ	Ã(_�NC�*��$�vA��p��ܸ�W�Du@C�IG��4��*I�m`�|�Ҙ<]�C�I<A��$#5厇M� Br	�?�VC�5"IB����V%����G�$i
C�I�+dTHI�Ǆ0n�����o��B�^��5���EdU��.�a��B�I�JD��)����GZ������B�I;� q�� �0.#,9[��\��C䉇SD��# �ҜoZ����"V��C�I$J��p�h�|i.�>br�C䉺:�x���n�O��	R��� zAjC�	�~� ����d�r�#ܐ>�&C�
UP���P�-<Ť�Cׂ�1-?*C�ɮ�9+������b���	�'��J�MAR*h�;�'��d�@8��'��#��T;I����eJ��0��'$Vٱ���!|��QV��x�H��'�D(1�Ɓ�l\�4l�th¥0�'N�ZS���'���.A�lA�'I�8�d�!.m̉+f��.�z��'����E�J�`�ʕ�6��{�`��'k,Ѩ cW*j�D�Jv�"e�9y�'�L�BA�8��m9��U�7�.ux��� ��@��
}8���T5G]� �7"OBl���`*Y ��W�j��!��"O�) ��s.�cf
�bވE��"Op!�CL�7j�E���ԿWY�Au"O`�K�ꋥ1�\���kI>^d�$�"O�ȳ�:$���(�-��Y�� �"ON�OC���YHeb�u�4� �"Ó���ͪ&��	Vk�0+�i0"O�ta�m�#@��M�qe¢���+g"O��F�	�v��|���_)0��@�0"O���!/ ��Y�lE)�ڴ8f"O�@�W��Y��|;!D�e��y�"O�؛�f[���`Cs�Љk}h"O-*�c�k�XyR���dx�#F"O�T���:h�`̀�)��V�A�a"O4��s�@{��k����kF�ax�"Od�; �%Q��I*˜�gfƱ�s"Od1���A��蘶KF+$QNx��"O6���n
1+Ѝ��
�v0b  "O���&��8� H���O�N�L��"O�!�g-�,L;��C�G�H=�[�"O��Ɂ�Ʈn�`R�&G'+-�y��"O�x���k��9�/�".%�!"O�Lq�H�V6�܊�+Ǜ>���k5"OdT�aaF�?� ��A׶GM�\�B"Oz ��.�8?�8�p����hMk�"OQQ����Dz�D^"�ܙ�"Of��e��O'�qJ�䚞y$�QQ"OdP��!O� �,e��S=lo8ٓ�"O
dj��j'.1���G�p��"OLAA����ɻa��<?���"OrP�d�G9~����&J]�4��8A"O�\)�U8(lBQ��7!f�,5"O����:o�u ���&e`��"O�P��샶�b �d�Y�Pg�B"O�9����A|)Z����!]n��A"Ox�)�BP�	ˆ��C[7ZV��剱b|�9��"SE���4DZ�r�^`a �3�B�
�Ԍr�Ƒ�	�ܔ2j"g{�,�@Ek�$�"~Γֈ�C��w����?4`�8�ȓ`��0��.�\^���ꉐ�B��Ik�N����^1l�a{�"X:��Ki݌a���8�L����=	�HJ�ƀih�bx� �:U.�h�$�Ƙ@��1;�"O�p��섺v�N�4)V,���E���'�V�XQ�)�D�G��ŉ�fxN�8! #�*�bF�	��yb�V�4�Ȝ�$c��+�F��I�6#f�*M�J72�'�>��}&�\�e H	{�ܜ�f-�h��B�ɌJUl�Q�L_�	�0p�e6�r�������1 Hְ=V���v	I%AZ�c�6� $.O����(�G���8v�io
��$���#�� j��&՜D��'�.e\� �L��Ri�7?��c��g��| �mXFj�x�OY�D��G�re�S��	8�� [�'s���P�PBv%���;���wgK�ߨ�1e$7}b��cG�9}0�[�� S(��B�O(D����S,0l�ewjA/*�X� �-�O>�*���r���
ۓ}�"95��cY����CX�O�ه�I�`IPR������cW�U��ACc�;�D(D�d��F�3y��� � �B�����&ʓdl��f!�'tm�1#c�V�+1��s�ّk �̄ȓ:��- ��۞=�
	��������ȓh�q���]�,�EE�O�&$�ȓ_�|�K�@(QFn���c��i;�)�ȓ>X@�Qvc�b�:��U�ƕm@�͆��zPZ��?��B�'��:� �%���>�F��O� �!����t�d���L�Z�LD�FO��b�"˓]#X	���e�,,�(�e��>9p��-����b6�ՊP-J`X�0Jd��bЛE�T?!+��@���ꐬ>ɐ4�fMX�<Ib�(�cb�I�Ȟ@��O�I�R��֋�OTG��A�X�t�����T��9��l���y�M<j�Xu��$�L��౑�9�����)�wy�g��?0�b?O�l��Ō=���9g�U.,��O*eh�`$t|�0	N0I`c�l!�GF������+q&�`1�\�B����F���ay��D�7� )Bg�L���H::&� ���2c�`5�1��!�+9V2t��h�nx�Mb� �/�'����d$�
uU��@���)�:|)���6p���c�_�zB��o�.G�˪�JH�� 
a�1ɦ+�!p���-��*��L<��G�Z?P ��i��,�V���QKh<1���Y`����'y�x:�L� ys���������f� ����'�<@�8�ϊ}ݤ=hc�B&A�V��鉾o��!Ba�`}�`��Gx���G��}��-م��o��YQԧ8y%a~Ҫ@��H�4AC�j���$hT��<1�C�(�'h�<�jF�fBҽ#I�n�Z���J�<Q���o���ꅿUlڬa���K�I}�Ȝ	c��(�?-q҇�#olA	P���UgŸ&"D�h�Ҭ�9����M�8h��0K�å.ȴ�c Z��Z�l�8
��<�B퉶G�|ysv�ҁH`�)�p��`
���R�Je�=�P��>1�k�Qovi�SLƴ/�X�8�U�o��y�4>�`���׾=���k �C)u1��G�k��'�V,��C�9҄���U� PTBЕ0x�')���ٿK	�T��%Nhņ�/���X��G z�����R�PN8`�蛍�~��^�*�.�r�
WܧJ�N� 5�¨9ra��B	څ
T��iPtO�H��h�N<����5.�1ʅ�z��X)P���~2�/'y.�#�
A�'O���E`V}���v*A�cU�T�
˓=�f�K�m� ®�\�V�0 �A� @F�`u�]���CG�Ōe��+��)h��Q����U�(~�u'�`#gY�f]�@�FU����m�a��'#g�1Ó�-s��a��E֮SJp�ȓ����ˇ�죑F$|Z��H`����D��6�"��%� J�� y�'�� ��F &��J�Ȕ�K0���'3�,(  &~r���o�� ^5 @�A�Hx±g�J?���a
8`�3ړ�D0 *[WҭC� 40~���IZSعk��@t}� ��Ri4&	�P��4fٖR4r��o4EeZ����1>��O��B�9p�*�)qxc�<`�j)	p�	�']m;$��+F��S�NX�ƩH�Z�(R��y�C�3%��t�T�)�̤8Ѯ[��OT�q�"��d+�5b���NV<ThE{g��0L6j�yB(�ze��%�(����>k�*T8��t�z��ȁy�b�O<��o�@�g�	!)(a�R��^��	ࢡ%tO��3��$&H�O1�@Rq�	m�"��@��U8L4�Bc������
��>�"�_�����:#z�)�>L,愦OD��ǒ��)�Y���CBG���䌇N�)e�+tB�T��hؚ3����C�o$��q
˷Sd�-�!i�)6vyb�����l+��.�J�����S�'	hd1� �	�$i����(W	�̇�	�$����˅y��	�O�sfLM�Nܱ)3�4,�����$�FE>� �l(y�ݝ i]�0
T&w��O����իJ8�9
�'Q�,5��i
����Zg��>Q=n���z��;$o�5��H� b��i��'A�D��r����L>1���0|0)�%�G�:���gr(<A'(�!�xM���&���d�?O�$|@��֖%���D�;]Mn(�-�=%<�� �x�ȷ�,@� �C~�#86�1�ս{�L!ч)��yb�������lU�%q�B�ēۢxc�����S�'S[���l���CF��27'T��s\��6��x�r�3D
t �����>>�?�'�>m _"dYz�͛�C��R��A�<I �2l���t�ʺra����U�<ٓ��\��٣" �q'��	�'�~�<� ���Sɛ3r,"P��%$Oj���"O�AQ����]�R����LH2��)b"O�.��z�������L6Խ9�"O��;U����@gH^*g>�H
�"O`UK&a0f�,ia�Fԫ7�hB'"Oʼ0���9����4B�+4�l�HF"O��r��5� 0
2�Y��A�g"O>x��K�-S��Ր��S�-Ȼ18O6�"�oڍ�p>���~�]��M�kX敡!-e��@������TΓ>{ ��򦂀{�F�SQ� �/ѐ�ȓ#Ӗx{��\5g�b����-DX�>�V놐U��Ts��!ڧP�v�P���\d(��Ḳ@f��ȓ'��)�c^�!�TdhtN�#u���IRK0~8�%
J�8��Y�L�ҡ�!4)�(�k�����e+D�\� �B�C�jd��l��s��i5�h��D�hR�J��hߓ`[�T8 ��5R�D�/ջ�8���J��� �%���[�&M����P�i����
�y�/Hc7�y��ףT�tl��.����'Yd� ��%*����^�V�á�~*�EFa��3	?&.��p+�|�<!�%E*Q]2 �&P�0��K�OqQF�BU� �Mc���w��銋�	�<�E�4T�*�Iviޡ�Tc�O�d�<��+��j�2�0G��h�n`
��A ��鈦�S�`w���͆&r��;l8��=!�SI��q�vA�5sɄ��A��X��X#��H��̌m����T��M
� P6��(��Pcl�:մ�)@�'L��6�ȼ?>�%��l6#`��p��$̻����xzr�+6eX�oC�ʧ}���P���g��9��@B���ȓ-Kȡ���D E(�he���'�X���G�8:����Y��2b�
NAp��4�tC�I0@�`����	gj�C��4'+Z5Sd��[�dCjDN��~&�d(���0���*�0Lz���.%�RC�ɂ������/J����C�J�RHk�\B*�r��'tB��h�>��}��鏾	;�A�˓@�À!S�tʓ��8��H�kh�΍0X1�ȓoD$� ���Ha��J�%�X!�Y#�N���:'!��P��D�"���Oq��C�ɋ��(h��&���� b��rе!�d�9�>�� ����B:"�hac��* �̬�ȓk3^<�$<G�;�R�(si��gil6JZ�VM��2J�mѦ���.�kU`��NNz��U��UҘ(��GN�D�B,	�Z��A��k6Y�ȓ��4r�iɪG������7n3�q��'��i���V"�@$ �0cό<�ȓ\�@�X�rE@�	�|�9�ȓN��X)q�X�j�, �n�
�,̄ȓi�v����v��(I��� �ȓ(UDb���[Ƣ� j5/�R��ȓp^ʩ�թʈS�H� ��ʤg}�I��FI�n	/JB�J��'s �`�ȓ|����C�r��c���y���ȓ!��DXU-�#Y�2�C2H�k��Q��DiHa�@㏏.���+�_�^��w�^1�"�!'���&�Aɦ̅ȓ!�d,��*T�k���\�^�,��ȓJk@u0�*6�X�CC��HS���`)Beѡ���Rۻi?�}�ȓ;Z
�Zed�9֚(F��	�vԇȓv��A@7�M�HXFp m��#G�����	uN�#DM_�
d��ȓ|�\YT�)���A��m�LY�ȓ@�ȵا!���e�cF�(ʺ���'p�:ŭ�-{ ���(��u	�!�ȓ�r�&�na�AQ�K��qЎх��v���CƵ�����(F��Ȇ�S�? � z!�O�I|ͫ�_�^�v"O6t�!л��\�D��6T�@T(w"OZ�
��Ro���Fɤl�8ɪ"O=k��-:��2ͮg���e�	�[Q�V�
5����-`��}��|�f&_�ju�h[�¦Z
��}�%3Ʈ�P|DA�T�ܸ���ȓv�ֹ��)�Y���۔p���'r6�6aJ,\�h鲅��-9�.���'��I��ؔCV|yZ�.��0�U�	�'e,��̗�)�n�[dO�"a&qJ�'�v�!5%S�u�t� ú&DD�{�'�P����V�	X�`�!Ʉ$,>���'���ٖ`�aR�q�$� �J�r�9�'�� �g�Ư\�DIZdS
A?}�K�������SD3���.�L�j��U�q��\Ǜ�%�	:C@	�A�|��i�eE !J�о<#��3��-$��QF$P"�ēZI���iT��<(��I
�A`��d N'7DA��'���^�q8尉��R:Jl����DY �c����v5t���F]Q?��]�D���۟�#}ZF�ӔA��#��:G����aG,e���r�(�{$�πYt��O�Q>� �^�yfE3���=W��q���>� �)��-���-}��	�稩j�E_x� �,Ț���*Y���'/}��<�d 3��ə�?�,���R��,�ҀL��M�C��(�qp ����ç]ܵ�V@D�0��8�
6!mrq���+oF����æE�6���0|��&�8v��U����H��r#@�\m��kg*|n���\�*6 �'>�}�FC΁Z&�$��#l4����e�n5����As�9�V�(Y4u��Sq�0���J�E��D��Q9EDѕ'���ELFd�͟X�?q[�.���؀�茥	RX���>au�F�Ff.IH��x���Ԣcذ\�C��5��d1��F5E��-��8���QC�'�~���� r���6�=a�'�8����/^�><�U�W�7� �'T��V �Ρ�A�5��Dx�'!����=
���J�
�%��U��'���!����D�<�R@�"�����'�8�Z��7XBxX�@��XDCO��yR����P���a�e^��y�C.2���� ����e���y��^c�HL��Eܺk h��.��y��c�Fm��/^(#���4�Y�yҥ�-gx���ED�!馘�S�ɑ�y�.Q$��m�gM�'�ȕ�#l̂�y�Lߏ:�fXb6aXzB�ț�R��y� G+!�̉YүC�BD�\�K��y���7�"̩ǀK�>�ɦ��/�y�k�$�6Xcw� �<��E�T��y�i�%�~��O&�"�+���y��ߚ1Y0Hp!h�U�H�����y�-ݦ$&�p8Rꚴc0Yxf����y2Kb�u(ϵ����uhR��y�ۯn��l����ʵiefA��yB�v}� #�8}���Y��yr�6f�P�i �!�T�ڄ�܊�yr(�h�C�)�r��휨�y�-P_�:�xC�#�a�Sdۖ�yrc�_����b7q`����`ڋ�yB�Ȫ� �3/�~^=��9�y�w�����|���3`���y���dYf��O,@�$�Ǒ�y�-L&�(͹� ���´#/I��yb.9;[x���+��H����y%�x����
	%.�t�Z箖!�y"��(}ܙk�y�� �$���yB�����bw�$^2̣����y�')z6THF坱 ���g�A�y�@ɏ\Pn=H�ַ�ĝf���y
� :�#���M#��"�^�g��H��"Oh@�F8|a�0�7jP�	�d� f"O�]�p�A 
��0)RIߛoEu�f"O���S��ri>1��(�q[�"O�����)oڑ�`�۱>%���t"O�lم�ۘI�f5:���"l|� �"O"�3��R���R�I��]�b"Oݠ�*�$yȐ f��-CnȨrw"O
��� X�X��H�dd%��"O��z����u���C�#rC� �"O6�Z��W;M��Pã��8$���H�"Ov��'d�Sk�\*0�D����"O&�84�D� \��Y���E��p�7"O�1�V�/���S�T�$�b���"O0�{'��A�J�a�б}���	�"O�͐��^U��e����}N�0�"O�jb�דG�>p#�AŢl����&"ON�$�1M?��@@.@-%�h�P"O`����8��葀&��S	|��"O���v	��yA�B+Ae桉!"O~�C���ɖ4�Ώ ~a��:$"O � ׌�6Y���������|"Oh��OA�5&<����>T�c"OV�!`�8l�lLX���=J����"OEEf]�e��lr ĝ3���Є"Oj!��T��a���Z�6�h�S"O��Q�փR��}�C�ԩf�Z��R"O���$�$j�q��yg��2�"O�U�QGZ`Ȝ�BFJ�3k�lu��"O�ъD��/J�� ����].TI��'�����J�&���cZ.\4 8��{�����+캩`0�)ZQd��ȓP�&��3��1�J��W&��3D�ę��B�~T���
��B��0ɣ�5D�@A�X'�h��P;*B���f6D���BP�_�v,���#����E�0D�@@��ĳ;}���_C ��kV)<D�|���
�6�s���-l"��
9D������
7`Y��E�>wD|i�$D�@�N`^H�;��
����G�#D��[e���!� �'�H�sK49 #�;D�Ls�/�+ar��a�F49'�r�?D�@z"'�%x9���!k����QKq�>D�� �Y�q� �x��� h��K��.D��$R��]=-Ҽ���0D��P��,o �(5c�����0w�8D��X!o ۆ\x7g$i|V #��p�<�J�9u�Kd�e64�f�HE�<)�� �	���b�⁽iJl\��O@�<���,W���1J�ǈ Çn�a�<��	����	�G͋X8"THT�Z؟��`<�ag�l�!��� /����ȓU�����ӑJ�䉪�`�l��\�ȓ8E�+�n%@Q�q-M2l��b�� wJ��=��H�s�X�|)��.r�+D�U�j�Pz��ߌ%����ul�)�˔"�Q*�ꁉ%*���J���z@�ŖN�@�B�l0�$��t3���FX����ҥ�u@V1��Q  ��E��
F��!ZD��o����	|�nG�TS�G������Fʥ %*]��G��1��H�Lϖ���M�d����^-�'��|��a4�+�FԆ��.@1ס�5{��)v��S�? t����1+{���a��,N�K�"O6�!�6�8�(�'ACL��#"O8�����/�L�EhǪ-lXٵ"O�h	��~6��7HG�`�a��"OZ�!"���8c�8�@��S�$9�Şoe�%q�J�x8�&��/{��ȓ:N*4�$�_ǮQ�\�!m����Y 昫� �'�(��"�V�%O,��H��0bvk�T��9�	�/W�lExr�'VVT�IQC��,{�^E#g�.�O����<�3._+1�&$�]�fǴl���C�<iՈA�{������s�]
0*�E�<���"~��{da�p"P��r@�f�<IǏǺSYy(5 �@�$2��f�<I�&��u��`������U�|�<i�*�5m��r�^�~� ���/u�<	$I�>+���X�GɤI��-�c�GF�<����f���C'�����0���B�<1�bK�f����T �l���`~�<�wi �O,�m(1�{X%�!�{�<�U�""��J�o�4y�"�X�����G{��	�0k�� Fn�90tev��p�C�ɩ(�sJ�U��Pe�HO.B�>���t*���T�pW�Ui�B��';O��ېE�t"�����<|�B�I�|�PhF.�}ช& ��8��B�ɐWH�P;�nB</�Ƽs�O?^f�B�Iwq��9!�ߦsJ�0�r�N��2C�I"c�cvB� �b�Q���r��C�	�H���"яf��YgO+)ۤC�ɴE��ɕd׆<ͬ�Ib̳S�C�ɪq�F�[�@W�FQ�%m��d�&C�I";��d�U'#k ��$dӶC�	�4|����LQ�#&ů	zC�	�m=r(9��4҈�G	E&2�B��n�������~ � �UB��<B�I?�p�ڀ�]ވ��iJ�H��B�� P���(EN�'ڠ�+VgE�~�B�I�]��(�+��,�� )V���B�I&8%z幅�_\����#��3��C�ɔ��ջ7A�R�.���
(j�*B�8r�d H3$�aC�ˆ�)��C�	�,�I:��D�F�y#���(��C�&K}4���⋌r����O�h��B�I%Z(@�%(� ��	�C�=��B�I@�*iI
�uD��ᔂ�(R�B䉑���wʷm;�aj0��.S�VC�I�@Lc#�K�Q±�cEE�<�C�ɩ{X�hS7��9=��֪�|��C䉨1��t� m��di���>C�	�d8�)�� ��S=Z|A�ʁ�*d(C�=4>&�i�j��zQ��"-�PB�	��*P�s��8�j���(U%\C䉆Qjl1E�"L4�5�["PO8C��
=�!�-F�-����B�	5�4X$�S=���Bj(&��C䉥H������ID�B��uGY,~޸B䉀?+)#thT� ��A�˖ZA�C�	n^��0S!Ég�آB�۶"Oz�%a���� 4��t��ta�"O0�HJ�3�Ā�UN��*b)��"O8�#�K���J=x n�"O!�$HM�
t��\?ϰ���gD0!�$� 'b�=�4$�2��Y�sH�q!�� .���)S��\�6�S�E 6���"O8 ��/�5w,�2����ѓ"O*��4F�?z�����	�g�ti�"O���`%��jHӓ��q�h��'"O�l�Po� a��h@��;3$�"T"Ol
A�S5�4؇M�:f+x]�"O���sf�m�QzPlK�G �M�t"On��S���ji��Sl�&hl�4"O��ӷ�/#�6,�'�0�u"O�3�铢n����	��X��"OD��5MF��Iy��4qU$83"O�,��ϋ��(P�����E��{"O�	"�Յ1��h��+'>f!{�"O��PB���\��(��'#�L(�"O@,�U�]!v�,I�V��)�)�P"O䭛cFB�\�I�`��1!�"�"O^1"���6I|�10Sc��Q&e�w"O�4b�Ȇ�D��x0�A�� �X)�a"O�]�"nĭc0eȤ��Z
�P��"OL��SmG�IdXpR�i�*q��"O�Z!E�?��+c��n��%"O���6e� =u����E���ԉ"O���4��R8�:�*$	~�`5"O��I�J��6����ޜ:AP�4"O81��Ɍ��JmR
Uv-�=rs"O&��D��q%�Y�G��	d-(4�c"O�����_,�N1#��0LE��"O�D�؉8\T�;�lA����Z�"O��Q�h��:�ΡK�@5`�ly%"O
U)D!Ʀ9��82#� ��j�"O��aC]"B�u9�\&�Dm�V"O��S��	��X$-W�4YuiF"O�@2h�1z�J� �Ҹ5!h����0��`�F��D芰L�A�p��6 ;�]Bce���(Od��J |s���A@M-9_��#�[�$�|����[�N�B-rc��wSͻ���>��O���DlU�s/h�*��1�(Uq�ؼD�^�6Gۅ9��]k�D�(+^�`��.Q�`�%��O�ąV�)̉Q\t�A�!�!����.*��	4>"\'���'����j�II�{R�s�,J<�̋E�'�7M~��E��T��S��>u���i�؟�z�46Q"��'^�L�'���A}��M������B:]8��܉���ۙ�tҴ�^��1#[�����-7q���ƫ0� �Ӡ�F [��C\���D�B[�L���S+!����R��Yt2�ydD�-~��*��}�㞉k�P�� v�X�0U�XӅ��O���TǦu�	H��6B#��<P��`��gD ���:wiV94��ٟ$������"�p�f���� w�J.Ց��mZ=�M���s�6�'���]qx���H�'h�UP��4/n����By�\�\Ҭ6M.�#�~Q۰G�N�e2�
�������.9
�@�gئI�Py`ՎVV��'
��c�D2D/#^B��,ӉR"��f��<C�ꕓ�C��
���"�w:r��C�K�D���0O���� �H2o�Z��`�;&�s���?����?�S�Y��⦝�&Ɛ1d����k�'w�v8:6�������Q��`z��#A�&M��!��&{�ꓩMS���������P{F�(��W�7ޔA��W`F�I�REɦ����T�� e,}�ᤇ�(�<��S$Ǡʓ��/<�H���D#���+��Ɏ%���"�����p7 	Լ�sf*5J�t����CjLT�r�"P���$�*�S��Ulڷ_Z"�
=���$\=7b�C��[ş���4�?�/Op��<�O|zAM�
�F�x&�7�N�p�l�I�<��`��` D	��S�ʈ0G*�~���ɦ�"۴��DJ�>�,�l�蟘�'$�T2w��k:��E�Z
N���D�O�[dk�*���<'Z�Ł>D�pt�e��:7`��S9�� i����d�"-1�O�\�Z��v�I8�p��M��sEd��%�.��!P�z�)i�ɢ%M"�D�O
Ql����;H�&	�7�>B<�UB�XL���?1)ON�S�O��ɢDXrж���-$��h���M��&˟|����JPo���8�DR-r�1,O��;�즅��~����R��p`QFI3}:���NK �I7R`1�ŉ�\Թ�w"�'ߘ�`���wX�MH�&N�
N��T'�ĄLr�Ox�iე�	���)�B������Þ(�U�P��� �����5Iۀ@�u�OvuV�L�d�O���S覝�	w�O��qS OM�RZ@��cj�ko�Y�I� ��N؞(�Q��Q�!�6*[�l��m���hOL4lZ�� $�$�;O�2��n�bu^XG�T/=&T�t�'k�'ay�%�5G $  �